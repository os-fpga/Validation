`include "encoder.v"
`include "invertion.v"
`include "large_adder.v"
`include "large_mux.v"
`include "memory_cntrl.v"
`include "register.v"
`include "full_adder.v"
`include "d_latch.v"
`include "shift_reg.v"
`include "mod_n_counter.v"
`include "decoder.v"
`include "parity_generator.v"

module design207_60_80_top #(parameter WIDTH=32,CHANNEL=60) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	reg [WIDTH-1:0] d_in10;
	reg [WIDTH-1:0] d_in11;
	reg [WIDTH-1:0] d_in12;
	reg [WIDTH-1:0] d_in13;
	reg [WIDTH-1:0] d_in14;
	reg [WIDTH-1:0] d_in15;
	reg [WIDTH-1:0] d_in16;
	reg [WIDTH-1:0] d_in17;
	reg [WIDTH-1:0] d_in18;
	reg [WIDTH-1:0] d_in19;
	reg [WIDTH-1:0] d_in20;
	reg [WIDTH-1:0] d_in21;
	reg [WIDTH-1:0] d_in22;
	reg [WIDTH-1:0] d_in23;
	reg [WIDTH-1:0] d_in24;
	reg [WIDTH-1:0] d_in25;
	reg [WIDTH-1:0] d_in26;
	reg [WIDTH-1:0] d_in27;
	reg [WIDTH-1:0] d_in28;
	reg [WIDTH-1:0] d_in29;
	reg [WIDTH-1:0] d_in30;
	reg [WIDTH-1:0] d_in31;
	reg [WIDTH-1:0] d_in32;
	reg [WIDTH-1:0] d_in33;
	reg [WIDTH-1:0] d_in34;
	reg [WIDTH-1:0] d_in35;
	reg [WIDTH-1:0] d_in36;
	reg [WIDTH-1:0] d_in37;
	reg [WIDTH-1:0] d_in38;
	reg [WIDTH-1:0] d_in39;
	reg [WIDTH-1:0] d_in40;
	reg [WIDTH-1:0] d_in41;
	reg [WIDTH-1:0] d_in42;
	reg [WIDTH-1:0] d_in43;
	reg [WIDTH-1:0] d_in44;
	reg [WIDTH-1:0] d_in45;
	reg [WIDTH-1:0] d_in46;
	reg [WIDTH-1:0] d_in47;
	reg [WIDTH-1:0] d_in48;
	reg [WIDTH-1:0] d_in49;
	reg [WIDTH-1:0] d_in50;
	reg [WIDTH-1:0] d_in51;
	reg [WIDTH-1:0] d_in52;
	reg [WIDTH-1:0] d_in53;
	reg [WIDTH-1:0] d_in54;
	reg [WIDTH-1:0] d_in55;
	reg [WIDTH-1:0] d_in56;
	reg [WIDTH-1:0] d_in57;
	reg [WIDTH-1:0] d_in58;
	reg [WIDTH-1:0] d_in59;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;
	wire [WIDTH-1:0] d_out10;
	wire [WIDTH-1:0] d_out11;
	wire [WIDTH-1:0] d_out12;
	wire [WIDTH-1:0] d_out13;
	wire [WIDTH-1:0] d_out14;
	wire [WIDTH-1:0] d_out15;
	wire [WIDTH-1:0] d_out16;
	wire [WIDTH-1:0] d_out17;
	wire [WIDTH-1:0] d_out18;
	wire [WIDTH-1:0] d_out19;
	wire [WIDTH-1:0] d_out20;
	wire [WIDTH-1:0] d_out21;
	wire [WIDTH-1:0] d_out22;
	wire [WIDTH-1:0] d_out23;
	wire [WIDTH-1:0] d_out24;
	wire [WIDTH-1:0] d_out25;
	wire [WIDTH-1:0] d_out26;
	wire [WIDTH-1:0] d_out27;
	wire [WIDTH-1:0] d_out28;
	wire [WIDTH-1:0] d_out29;
	wire [WIDTH-1:0] d_out30;
	wire [WIDTH-1:0] d_out31;
	wire [WIDTH-1:0] d_out32;
	wire [WIDTH-1:0] d_out33;
	wire [WIDTH-1:0] d_out34;
	wire [WIDTH-1:0] d_out35;
	wire [WIDTH-1:0] d_out36;
	wire [WIDTH-1:0] d_out37;
	wire [WIDTH-1:0] d_out38;
	wire [WIDTH-1:0] d_out39;
	wire [WIDTH-1:0] d_out40;
	wire [WIDTH-1:0] d_out41;
	wire [WIDTH-1:0] d_out42;
	wire [WIDTH-1:0] d_out43;
	wire [WIDTH-1:0] d_out44;
	wire [WIDTH-1:0] d_out45;
	wire [WIDTH-1:0] d_out46;
	wire [WIDTH-1:0] d_out47;
	wire [WIDTH-1:0] d_out48;
	wire [WIDTH-1:0] d_out49;
	wire [WIDTH-1:0] d_out50;
	wire [WIDTH-1:0] d_out51;
	wire [WIDTH-1:0] d_out52;
	wire [WIDTH-1:0] d_out53;
	wire [WIDTH-1:0] d_out54;
	wire [WIDTH-1:0] d_out55;
	wire [WIDTH-1:0] d_out56;
	wire [WIDTH-1:0] d_out57;
	wire [WIDTH-1:0] d_out58;
	wire [WIDTH-1:0] d_out59;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH-1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 <= tmp[WIDTH-1:0];
		d_in1 <= tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 <= tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 <= tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 <= tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 <= tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 <= tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 <= tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 <= tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 <= tmp[(WIDTH*10)-1:WIDTH*9];
		d_in10 <= tmp[(WIDTH*11)-1:WIDTH*10];
		d_in11 <= tmp[(WIDTH*12)-1:WIDTH*11];
		d_in12 <= tmp[(WIDTH*13)-1:WIDTH*12];
		d_in13 <= tmp[(WIDTH*14)-1:WIDTH*13];
		d_in14 <= tmp[(WIDTH*15)-1:WIDTH*14];
		d_in15 <= tmp[(WIDTH*16)-1:WIDTH*15];
		d_in16 <= tmp[(WIDTH*17)-1:WIDTH*16];
		d_in17 <= tmp[(WIDTH*18)-1:WIDTH*17];
		d_in18 <= tmp[(WIDTH*19)-1:WIDTH*18];
		d_in19 <= tmp[(WIDTH*20)-1:WIDTH*19];
		d_in20 <= tmp[(WIDTH*21)-1:WIDTH*20];
		d_in21 <= tmp[(WIDTH*22)-1:WIDTH*21];
		d_in22 <= tmp[(WIDTH*23)-1:WIDTH*22];
		d_in23 <= tmp[(WIDTH*24)-1:WIDTH*23];
		d_in24 <= tmp[(WIDTH*25)-1:WIDTH*24];
		d_in25 <= tmp[(WIDTH*26)-1:WIDTH*25];
		d_in26 <= tmp[(WIDTH*27)-1:WIDTH*26];
		d_in27 <= tmp[(WIDTH*28)-1:WIDTH*27];
		d_in28 <= tmp[(WIDTH*29)-1:WIDTH*28];
		d_in29 <= tmp[(WIDTH*30)-1:WIDTH*29];
		d_in30 <= tmp[(WIDTH*31)-1:WIDTH*30];
		d_in31 <= tmp[(WIDTH*32)-1:WIDTH*31];
		d_in32 <= tmp[(WIDTH*33)-1:WIDTH*32];
		d_in33 <= tmp[(WIDTH*34)-1:WIDTH*33];
		d_in34 <= tmp[(WIDTH*35)-1:WIDTH*34];
		d_in35 <= tmp[(WIDTH*36)-1:WIDTH*35];
		d_in36 <= tmp[(WIDTH*37)-1:WIDTH*36];
		d_in37 <= tmp[(WIDTH*38)-1:WIDTH*37];
		d_in38 <= tmp[(WIDTH*39)-1:WIDTH*38];
		d_in39 <= tmp[(WIDTH*40)-1:WIDTH*39];
		d_in40 <= tmp[(WIDTH*41)-1:WIDTH*40];
		d_in41 <= tmp[(WIDTH*42)-1:WIDTH*41];
		d_in42 <= tmp[(WIDTH*43)-1:WIDTH*42];
		d_in43 <= tmp[(WIDTH*44)-1:WIDTH*43];
		d_in44 <= tmp[(WIDTH*45)-1:WIDTH*44];
		d_in45 <= tmp[(WIDTH*46)-1:WIDTH*45];
		d_in46 <= tmp[(WIDTH*47)-1:WIDTH*46];
		d_in47 <= tmp[(WIDTH*48)-1:WIDTH*47];
		d_in48 <= tmp[(WIDTH*49)-1:WIDTH*48];
		d_in49 <= tmp[(WIDTH*50)-1:WIDTH*49];
		d_in50 <= tmp[(WIDTH*51)-1:WIDTH*50];
		d_in51 <= tmp[(WIDTH*52)-1:WIDTH*51];
		d_in52 <= tmp[(WIDTH*53)-1:WIDTH*52];
		d_in53 <= tmp[(WIDTH*54)-1:WIDTH*53];
		d_in54 <= tmp[(WIDTH*55)-1:WIDTH*54];
		d_in55 <= tmp[(WIDTH*56)-1:WIDTH*55];
		d_in56 <= tmp[(WIDTH*57)-1:WIDTH*56];
		d_in57 <= tmp[(WIDTH*58)-1:WIDTH*57];
		d_in58 <= tmp[(WIDTH*59)-1:WIDTH*58];
		d_in59 <= tmp[(WIDTH*60)-1:WIDTH*59];
	end

	design207_60_80 #(.WIDTH(WIDTH)) design207_60_80_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_in10(d_in10),.d_in11(d_in11),.d_in12(d_in12),.d_in13(d_in13),.d_in14(d_in14),.d_in15(d_in15),.d_in16(d_in16),.d_in17(d_in17),.d_in18(d_in18),.d_in19(d_in19),.d_in20(d_in20),.d_in21(d_in21),.d_in22(d_in22),.d_in23(d_in23),.d_in24(d_in24),.d_in25(d_in25),.d_in26(d_in26),.d_in27(d_in27),.d_in28(d_in28),.d_in29(d_in29),.d_in30(d_in30),.d_in31(d_in31),.d_in32(d_in32),.d_in33(d_in33),.d_in34(d_in34),.d_in35(d_in35),.d_in36(d_in36),.d_in37(d_in37),.d_in38(d_in38),.d_in39(d_in39),.d_in40(d_in40),.d_in41(d_in41),.d_in42(d_in42),.d_in43(d_in43),.d_in44(d_in44),.d_in45(d_in45),.d_in46(d_in46),.d_in47(d_in47),.d_in48(d_in48),.d_in49(d_in49),.d_in50(d_in50),.d_in51(d_in51),.d_in52(d_in52),.d_in53(d_in53),.d_in54(d_in54),.d_in55(d_in55),.d_in56(d_in56),.d_in57(d_in57),.d_in58(d_in58),.d_in59(d_in59),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.d_out10(d_out10),.d_out11(d_out11),.d_out12(d_out12),.d_out13(d_out13),.d_out14(d_out14),.d_out15(d_out15),.d_out16(d_out16),.d_out17(d_out17),.d_out18(d_out18),.d_out19(d_out19),.d_out20(d_out20),.d_out21(d_out21),.d_out22(d_out22),.d_out23(d_out23),.d_out24(d_out24),.d_out25(d_out25),.d_out26(d_out26),.d_out27(d_out27),.d_out28(d_out28),.d_out29(d_out29),.d_out30(d_out30),.d_out31(d_out31),.d_out32(d_out32),.d_out33(d_out33),.d_out34(d_out34),.d_out35(d_out35),.d_out36(d_out36),.d_out37(d_out37),.d_out38(d_out38),.d_out39(d_out39),.d_out40(d_out40),.d_out41(d_out41),.d_out42(d_out42),.d_out43(d_out43),.d_out44(d_out44),.d_out45(d_out45),.d_out46(d_out46),.d_out47(d_out47),.d_out48(d_out48),.d_out49(d_out49),.d_out50(d_out50),.d_out51(d_out51),.d_out52(d_out52),.d_out53(d_out53),.d_out54(d_out54),.d_out55(d_out55),.d_out56(d_out56),.d_out57(d_out57),.d_out58(d_out58),.d_out59(d_out59),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9^d_out10^d_out11^d_out12^d_out13^d_out14^d_out15^d_out16^d_out17^d_out18^d_out19^d_out20^d_out21^d_out22^d_out23^d_out24^d_out25^d_out26^d_out27^d_out28^d_out29^d_out30^d_out31^d_out32^d_out33^d_out34^d_out35^d_out36^d_out37^d_out38^d_out39^d_out40^d_out41^d_out42^d_out43^d_out44^d_out45^d_out46^d_out47^d_out48^d_out49^d_out50^d_out51^d_out52^d_out53^d_out54^d_out55^d_out56^d_out57^d_out58^d_out59;

endmodule

module design207_60_80 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_in10, d_in11, d_in12, d_in13, d_in14, d_in15, d_in16, d_in17, d_in18, d_in19, d_in20, d_in21, d_in22, d_in23, d_in24, d_in25, d_in26, d_in27, d_in28, d_in29, d_in30, d_in31, d_in32, d_in33, d_in34, d_in35, d_in36, d_in37, d_in38, d_in39, d_in40, d_in41, d_in42, d_in43, d_in44, d_in45, d_in46, d_in47, d_in48, d_in49, d_in50, d_in51, d_in52, d_in53, d_in54, d_in55, d_in56, d_in57, d_in58, d_in59, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, d_out10, d_out11, d_out12, d_out13, d_out14, d_out15, d_out16, d_out17, d_out18, d_out19, d_out20, d_out21, d_out22, d_out23, d_out24, d_out25, d_out26, d_out27, d_out28, d_out29, d_out30, d_out31, d_out32, d_out33, d_out34, d_out35, d_out36, d_out37, d_out38, d_out39, d_out40, d_out41, d_out42, d_out43, d_out44, d_out45, d_out46, d_out47, d_out48, d_out49, d_out50, d_out51, d_out52, d_out53, d_out54, d_out55, d_out56, d_out57, d_out58, d_out59, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	input [WIDTH-1:0] d_in10; 
	input [WIDTH-1:0] d_in11; 
	input [WIDTH-1:0] d_in12; 
	input [WIDTH-1:0] d_in13; 
	input [WIDTH-1:0] d_in14; 
	input [WIDTH-1:0] d_in15; 
	input [WIDTH-1:0] d_in16; 
	input [WIDTH-1:0] d_in17; 
	input [WIDTH-1:0] d_in18; 
	input [WIDTH-1:0] d_in19; 
	input [WIDTH-1:0] d_in20; 
	input [WIDTH-1:0] d_in21; 
	input [WIDTH-1:0] d_in22; 
	input [WIDTH-1:0] d_in23; 
	input [WIDTH-1:0] d_in24; 
	input [WIDTH-1:0] d_in25; 
	input [WIDTH-1:0] d_in26; 
	input [WIDTH-1:0] d_in27; 
	input [WIDTH-1:0] d_in28; 
	input [WIDTH-1:0] d_in29; 
	input [WIDTH-1:0] d_in30; 
	input [WIDTH-1:0] d_in31; 
	input [WIDTH-1:0] d_in32; 
	input [WIDTH-1:0] d_in33; 
	input [WIDTH-1:0] d_in34; 
	input [WIDTH-1:0] d_in35; 
	input [WIDTH-1:0] d_in36; 
	input [WIDTH-1:0] d_in37; 
	input [WIDTH-1:0] d_in38; 
	input [WIDTH-1:0] d_in39; 
	input [WIDTH-1:0] d_in40; 
	input [WIDTH-1:0] d_in41; 
	input [WIDTH-1:0] d_in42; 
	input [WIDTH-1:0] d_in43; 
	input [WIDTH-1:0] d_in44; 
	input [WIDTH-1:0] d_in45; 
	input [WIDTH-1:0] d_in46; 
	input [WIDTH-1:0] d_in47; 
	input [WIDTH-1:0] d_in48; 
	input [WIDTH-1:0] d_in49; 
	input [WIDTH-1:0] d_in50; 
	input [WIDTH-1:0] d_in51; 
	input [WIDTH-1:0] d_in52; 
	input [WIDTH-1:0] d_in53; 
	input [WIDTH-1:0] d_in54; 
	input [WIDTH-1:0] d_in55; 
	input [WIDTH-1:0] d_in56; 
	input [WIDTH-1:0] d_in57; 
	input [WIDTH-1:0] d_in58; 
	input [WIDTH-1:0] d_in59; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 
	output [WIDTH-1:0] d_out10; 
	output [WIDTH-1:0] d_out11; 
	output [WIDTH-1:0] d_out12; 
	output [WIDTH-1:0] d_out13; 
	output [WIDTH-1:0] d_out14; 
	output [WIDTH-1:0] d_out15; 
	output [WIDTH-1:0] d_out16; 
	output [WIDTH-1:0] d_out17; 
	output [WIDTH-1:0] d_out18; 
	output [WIDTH-1:0] d_out19; 
	output [WIDTH-1:0] d_out20; 
	output [WIDTH-1:0] d_out21; 
	output [WIDTH-1:0] d_out22; 
	output [WIDTH-1:0] d_out23; 
	output [WIDTH-1:0] d_out24; 
	output [WIDTH-1:0] d_out25; 
	output [WIDTH-1:0] d_out26; 
	output [WIDTH-1:0] d_out27; 
	output [WIDTH-1:0] d_out28; 
	output [WIDTH-1:0] d_out29; 
	output [WIDTH-1:0] d_out30; 
	output [WIDTH-1:0] d_out31; 
	output [WIDTH-1:0] d_out32; 
	output [WIDTH-1:0] d_out33; 
	output [WIDTH-1:0] d_out34; 
	output [WIDTH-1:0] d_out35; 
	output [WIDTH-1:0] d_out36; 
	output [WIDTH-1:0] d_out37; 
	output [WIDTH-1:0] d_out38; 
	output [WIDTH-1:0] d_out39; 
	output [WIDTH-1:0] d_out40; 
	output [WIDTH-1:0] d_out41; 
	output [WIDTH-1:0] d_out42; 
	output [WIDTH-1:0] d_out43; 
	output [WIDTH-1:0] d_out44; 
	output [WIDTH-1:0] d_out45; 
	output [WIDTH-1:0] d_out46; 
	output [WIDTH-1:0] d_out47; 
	output [WIDTH-1:0] d_out48; 
	output [WIDTH-1:0] d_out49; 
	output [WIDTH-1:0] d_out50; 
	output [WIDTH-1:0] d_out51; 
	output [WIDTH-1:0] d_out52; 
	output [WIDTH-1:0] d_out53; 
	output [WIDTH-1:0] d_out54; 
	output [WIDTH-1:0] d_out55; 
	output [WIDTH-1:0] d_out56; 
	output [WIDTH-1:0] d_out57; 
	output [WIDTH-1:0] d_out58; 
	output [WIDTH-1:0] d_out59; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d0_29;
	wire [WIDTH-1:0] wire_d0_30;
	wire [WIDTH-1:0] wire_d0_31;
	wire [WIDTH-1:0] wire_d0_32;
	wire [WIDTH-1:0] wire_d0_33;
	wire [WIDTH-1:0] wire_d0_34;
	wire [WIDTH-1:0] wire_d0_35;
	wire [WIDTH-1:0] wire_d0_36;
	wire [WIDTH-1:0] wire_d0_37;
	wire [WIDTH-1:0] wire_d0_38;
	wire [WIDTH-1:0] wire_d0_39;
	wire [WIDTH-1:0] wire_d0_40;
	wire [WIDTH-1:0] wire_d0_41;
	wire [WIDTH-1:0] wire_d0_42;
	wire [WIDTH-1:0] wire_d0_43;
	wire [WIDTH-1:0] wire_d0_44;
	wire [WIDTH-1:0] wire_d0_45;
	wire [WIDTH-1:0] wire_d0_46;
	wire [WIDTH-1:0] wire_d0_47;
	wire [WIDTH-1:0] wire_d0_48;
	wire [WIDTH-1:0] wire_d0_49;
	wire [WIDTH-1:0] wire_d0_50;
	wire [WIDTH-1:0] wire_d0_51;
	wire [WIDTH-1:0] wire_d0_52;
	wire [WIDTH-1:0] wire_d0_53;
	wire [WIDTH-1:0] wire_d0_54;
	wire [WIDTH-1:0] wire_d0_55;
	wire [WIDTH-1:0] wire_d0_56;
	wire [WIDTH-1:0] wire_d0_57;
	wire [WIDTH-1:0] wire_d0_58;
	wire [WIDTH-1:0] wire_d0_59;
	wire [WIDTH-1:0] wire_d0_60;
	wire [WIDTH-1:0] wire_d0_61;
	wire [WIDTH-1:0] wire_d0_62;
	wire [WIDTH-1:0] wire_d0_63;
	wire [WIDTH-1:0] wire_d0_64;
	wire [WIDTH-1:0] wire_d0_65;
	wire [WIDTH-1:0] wire_d0_66;
	wire [WIDTH-1:0] wire_d0_67;
	wire [WIDTH-1:0] wire_d0_68;
	wire [WIDTH-1:0] wire_d0_69;
	wire [WIDTH-1:0] wire_d0_70;
	wire [WIDTH-1:0] wire_d0_71;
	wire [WIDTH-1:0] wire_d0_72;
	wire [WIDTH-1:0] wire_d0_73;
	wire [WIDTH-1:0] wire_d0_74;
	wire [WIDTH-1:0] wire_d0_75;
	wire [WIDTH-1:0] wire_d0_76;
	wire [WIDTH-1:0] wire_d0_77;
	wire [WIDTH-1:0] wire_d0_78;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d1_29;
	wire [WIDTH-1:0] wire_d1_30;
	wire [WIDTH-1:0] wire_d1_31;
	wire [WIDTH-1:0] wire_d1_32;
	wire [WIDTH-1:0] wire_d1_33;
	wire [WIDTH-1:0] wire_d1_34;
	wire [WIDTH-1:0] wire_d1_35;
	wire [WIDTH-1:0] wire_d1_36;
	wire [WIDTH-1:0] wire_d1_37;
	wire [WIDTH-1:0] wire_d1_38;
	wire [WIDTH-1:0] wire_d1_39;
	wire [WIDTH-1:0] wire_d1_40;
	wire [WIDTH-1:0] wire_d1_41;
	wire [WIDTH-1:0] wire_d1_42;
	wire [WIDTH-1:0] wire_d1_43;
	wire [WIDTH-1:0] wire_d1_44;
	wire [WIDTH-1:0] wire_d1_45;
	wire [WIDTH-1:0] wire_d1_46;
	wire [WIDTH-1:0] wire_d1_47;
	wire [WIDTH-1:0] wire_d1_48;
	wire [WIDTH-1:0] wire_d1_49;
	wire [WIDTH-1:0] wire_d1_50;
	wire [WIDTH-1:0] wire_d1_51;
	wire [WIDTH-1:0] wire_d1_52;
	wire [WIDTH-1:0] wire_d1_53;
	wire [WIDTH-1:0] wire_d1_54;
	wire [WIDTH-1:0] wire_d1_55;
	wire [WIDTH-1:0] wire_d1_56;
	wire [WIDTH-1:0] wire_d1_57;
	wire [WIDTH-1:0] wire_d1_58;
	wire [WIDTH-1:0] wire_d1_59;
	wire [WIDTH-1:0] wire_d1_60;
	wire [WIDTH-1:0] wire_d1_61;
	wire [WIDTH-1:0] wire_d1_62;
	wire [WIDTH-1:0] wire_d1_63;
	wire [WIDTH-1:0] wire_d1_64;
	wire [WIDTH-1:0] wire_d1_65;
	wire [WIDTH-1:0] wire_d1_66;
	wire [WIDTH-1:0] wire_d1_67;
	wire [WIDTH-1:0] wire_d1_68;
	wire [WIDTH-1:0] wire_d1_69;
	wire [WIDTH-1:0] wire_d1_70;
	wire [WIDTH-1:0] wire_d1_71;
	wire [WIDTH-1:0] wire_d1_72;
	wire [WIDTH-1:0] wire_d1_73;
	wire [WIDTH-1:0] wire_d1_74;
	wire [WIDTH-1:0] wire_d1_75;
	wire [WIDTH-1:0] wire_d1_76;
	wire [WIDTH-1:0] wire_d1_77;
	wire [WIDTH-1:0] wire_d1_78;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d2_29;
	wire [WIDTH-1:0] wire_d2_30;
	wire [WIDTH-1:0] wire_d2_31;
	wire [WIDTH-1:0] wire_d2_32;
	wire [WIDTH-1:0] wire_d2_33;
	wire [WIDTH-1:0] wire_d2_34;
	wire [WIDTH-1:0] wire_d2_35;
	wire [WIDTH-1:0] wire_d2_36;
	wire [WIDTH-1:0] wire_d2_37;
	wire [WIDTH-1:0] wire_d2_38;
	wire [WIDTH-1:0] wire_d2_39;
	wire [WIDTH-1:0] wire_d2_40;
	wire [WIDTH-1:0] wire_d2_41;
	wire [WIDTH-1:0] wire_d2_42;
	wire [WIDTH-1:0] wire_d2_43;
	wire [WIDTH-1:0] wire_d2_44;
	wire [WIDTH-1:0] wire_d2_45;
	wire [WIDTH-1:0] wire_d2_46;
	wire [WIDTH-1:0] wire_d2_47;
	wire [WIDTH-1:0] wire_d2_48;
	wire [WIDTH-1:0] wire_d2_49;
	wire [WIDTH-1:0] wire_d2_50;
	wire [WIDTH-1:0] wire_d2_51;
	wire [WIDTH-1:0] wire_d2_52;
	wire [WIDTH-1:0] wire_d2_53;
	wire [WIDTH-1:0] wire_d2_54;
	wire [WIDTH-1:0] wire_d2_55;
	wire [WIDTH-1:0] wire_d2_56;
	wire [WIDTH-1:0] wire_d2_57;
	wire [WIDTH-1:0] wire_d2_58;
	wire [WIDTH-1:0] wire_d2_59;
	wire [WIDTH-1:0] wire_d2_60;
	wire [WIDTH-1:0] wire_d2_61;
	wire [WIDTH-1:0] wire_d2_62;
	wire [WIDTH-1:0] wire_d2_63;
	wire [WIDTH-1:0] wire_d2_64;
	wire [WIDTH-1:0] wire_d2_65;
	wire [WIDTH-1:0] wire_d2_66;
	wire [WIDTH-1:0] wire_d2_67;
	wire [WIDTH-1:0] wire_d2_68;
	wire [WIDTH-1:0] wire_d2_69;
	wire [WIDTH-1:0] wire_d2_70;
	wire [WIDTH-1:0] wire_d2_71;
	wire [WIDTH-1:0] wire_d2_72;
	wire [WIDTH-1:0] wire_d2_73;
	wire [WIDTH-1:0] wire_d2_74;
	wire [WIDTH-1:0] wire_d2_75;
	wire [WIDTH-1:0] wire_d2_76;
	wire [WIDTH-1:0] wire_d2_77;
	wire [WIDTH-1:0] wire_d2_78;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d3_29;
	wire [WIDTH-1:0] wire_d3_30;
	wire [WIDTH-1:0] wire_d3_31;
	wire [WIDTH-1:0] wire_d3_32;
	wire [WIDTH-1:0] wire_d3_33;
	wire [WIDTH-1:0] wire_d3_34;
	wire [WIDTH-1:0] wire_d3_35;
	wire [WIDTH-1:0] wire_d3_36;
	wire [WIDTH-1:0] wire_d3_37;
	wire [WIDTH-1:0] wire_d3_38;
	wire [WIDTH-1:0] wire_d3_39;
	wire [WIDTH-1:0] wire_d3_40;
	wire [WIDTH-1:0] wire_d3_41;
	wire [WIDTH-1:0] wire_d3_42;
	wire [WIDTH-1:0] wire_d3_43;
	wire [WIDTH-1:0] wire_d3_44;
	wire [WIDTH-1:0] wire_d3_45;
	wire [WIDTH-1:0] wire_d3_46;
	wire [WIDTH-1:0] wire_d3_47;
	wire [WIDTH-1:0] wire_d3_48;
	wire [WIDTH-1:0] wire_d3_49;
	wire [WIDTH-1:0] wire_d3_50;
	wire [WIDTH-1:0] wire_d3_51;
	wire [WIDTH-1:0] wire_d3_52;
	wire [WIDTH-1:0] wire_d3_53;
	wire [WIDTH-1:0] wire_d3_54;
	wire [WIDTH-1:0] wire_d3_55;
	wire [WIDTH-1:0] wire_d3_56;
	wire [WIDTH-1:0] wire_d3_57;
	wire [WIDTH-1:0] wire_d3_58;
	wire [WIDTH-1:0] wire_d3_59;
	wire [WIDTH-1:0] wire_d3_60;
	wire [WIDTH-1:0] wire_d3_61;
	wire [WIDTH-1:0] wire_d3_62;
	wire [WIDTH-1:0] wire_d3_63;
	wire [WIDTH-1:0] wire_d3_64;
	wire [WIDTH-1:0] wire_d3_65;
	wire [WIDTH-1:0] wire_d3_66;
	wire [WIDTH-1:0] wire_d3_67;
	wire [WIDTH-1:0] wire_d3_68;
	wire [WIDTH-1:0] wire_d3_69;
	wire [WIDTH-1:0] wire_d3_70;
	wire [WIDTH-1:0] wire_d3_71;
	wire [WIDTH-1:0] wire_d3_72;
	wire [WIDTH-1:0] wire_d3_73;
	wire [WIDTH-1:0] wire_d3_74;
	wire [WIDTH-1:0] wire_d3_75;
	wire [WIDTH-1:0] wire_d3_76;
	wire [WIDTH-1:0] wire_d3_77;
	wire [WIDTH-1:0] wire_d3_78;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d4_29;
	wire [WIDTH-1:0] wire_d4_30;
	wire [WIDTH-1:0] wire_d4_31;
	wire [WIDTH-1:0] wire_d4_32;
	wire [WIDTH-1:0] wire_d4_33;
	wire [WIDTH-1:0] wire_d4_34;
	wire [WIDTH-1:0] wire_d4_35;
	wire [WIDTH-1:0] wire_d4_36;
	wire [WIDTH-1:0] wire_d4_37;
	wire [WIDTH-1:0] wire_d4_38;
	wire [WIDTH-1:0] wire_d4_39;
	wire [WIDTH-1:0] wire_d4_40;
	wire [WIDTH-1:0] wire_d4_41;
	wire [WIDTH-1:0] wire_d4_42;
	wire [WIDTH-1:0] wire_d4_43;
	wire [WIDTH-1:0] wire_d4_44;
	wire [WIDTH-1:0] wire_d4_45;
	wire [WIDTH-1:0] wire_d4_46;
	wire [WIDTH-1:0] wire_d4_47;
	wire [WIDTH-1:0] wire_d4_48;
	wire [WIDTH-1:0] wire_d4_49;
	wire [WIDTH-1:0] wire_d4_50;
	wire [WIDTH-1:0] wire_d4_51;
	wire [WIDTH-1:0] wire_d4_52;
	wire [WIDTH-1:0] wire_d4_53;
	wire [WIDTH-1:0] wire_d4_54;
	wire [WIDTH-1:0] wire_d4_55;
	wire [WIDTH-1:0] wire_d4_56;
	wire [WIDTH-1:0] wire_d4_57;
	wire [WIDTH-1:0] wire_d4_58;
	wire [WIDTH-1:0] wire_d4_59;
	wire [WIDTH-1:0] wire_d4_60;
	wire [WIDTH-1:0] wire_d4_61;
	wire [WIDTH-1:0] wire_d4_62;
	wire [WIDTH-1:0] wire_d4_63;
	wire [WIDTH-1:0] wire_d4_64;
	wire [WIDTH-1:0] wire_d4_65;
	wire [WIDTH-1:0] wire_d4_66;
	wire [WIDTH-1:0] wire_d4_67;
	wire [WIDTH-1:0] wire_d4_68;
	wire [WIDTH-1:0] wire_d4_69;
	wire [WIDTH-1:0] wire_d4_70;
	wire [WIDTH-1:0] wire_d4_71;
	wire [WIDTH-1:0] wire_d4_72;
	wire [WIDTH-1:0] wire_d4_73;
	wire [WIDTH-1:0] wire_d4_74;
	wire [WIDTH-1:0] wire_d4_75;
	wire [WIDTH-1:0] wire_d4_76;
	wire [WIDTH-1:0] wire_d4_77;
	wire [WIDTH-1:0] wire_d4_78;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d5_29;
	wire [WIDTH-1:0] wire_d5_30;
	wire [WIDTH-1:0] wire_d5_31;
	wire [WIDTH-1:0] wire_d5_32;
	wire [WIDTH-1:0] wire_d5_33;
	wire [WIDTH-1:0] wire_d5_34;
	wire [WIDTH-1:0] wire_d5_35;
	wire [WIDTH-1:0] wire_d5_36;
	wire [WIDTH-1:0] wire_d5_37;
	wire [WIDTH-1:0] wire_d5_38;
	wire [WIDTH-1:0] wire_d5_39;
	wire [WIDTH-1:0] wire_d5_40;
	wire [WIDTH-1:0] wire_d5_41;
	wire [WIDTH-1:0] wire_d5_42;
	wire [WIDTH-1:0] wire_d5_43;
	wire [WIDTH-1:0] wire_d5_44;
	wire [WIDTH-1:0] wire_d5_45;
	wire [WIDTH-1:0] wire_d5_46;
	wire [WIDTH-1:0] wire_d5_47;
	wire [WIDTH-1:0] wire_d5_48;
	wire [WIDTH-1:0] wire_d5_49;
	wire [WIDTH-1:0] wire_d5_50;
	wire [WIDTH-1:0] wire_d5_51;
	wire [WIDTH-1:0] wire_d5_52;
	wire [WIDTH-1:0] wire_d5_53;
	wire [WIDTH-1:0] wire_d5_54;
	wire [WIDTH-1:0] wire_d5_55;
	wire [WIDTH-1:0] wire_d5_56;
	wire [WIDTH-1:0] wire_d5_57;
	wire [WIDTH-1:0] wire_d5_58;
	wire [WIDTH-1:0] wire_d5_59;
	wire [WIDTH-1:0] wire_d5_60;
	wire [WIDTH-1:0] wire_d5_61;
	wire [WIDTH-1:0] wire_d5_62;
	wire [WIDTH-1:0] wire_d5_63;
	wire [WIDTH-1:0] wire_d5_64;
	wire [WIDTH-1:0] wire_d5_65;
	wire [WIDTH-1:0] wire_d5_66;
	wire [WIDTH-1:0] wire_d5_67;
	wire [WIDTH-1:0] wire_d5_68;
	wire [WIDTH-1:0] wire_d5_69;
	wire [WIDTH-1:0] wire_d5_70;
	wire [WIDTH-1:0] wire_d5_71;
	wire [WIDTH-1:0] wire_d5_72;
	wire [WIDTH-1:0] wire_d5_73;
	wire [WIDTH-1:0] wire_d5_74;
	wire [WIDTH-1:0] wire_d5_75;
	wire [WIDTH-1:0] wire_d5_76;
	wire [WIDTH-1:0] wire_d5_77;
	wire [WIDTH-1:0] wire_d5_78;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d6_29;
	wire [WIDTH-1:0] wire_d6_30;
	wire [WIDTH-1:0] wire_d6_31;
	wire [WIDTH-1:0] wire_d6_32;
	wire [WIDTH-1:0] wire_d6_33;
	wire [WIDTH-1:0] wire_d6_34;
	wire [WIDTH-1:0] wire_d6_35;
	wire [WIDTH-1:0] wire_d6_36;
	wire [WIDTH-1:0] wire_d6_37;
	wire [WIDTH-1:0] wire_d6_38;
	wire [WIDTH-1:0] wire_d6_39;
	wire [WIDTH-1:0] wire_d6_40;
	wire [WIDTH-1:0] wire_d6_41;
	wire [WIDTH-1:0] wire_d6_42;
	wire [WIDTH-1:0] wire_d6_43;
	wire [WIDTH-1:0] wire_d6_44;
	wire [WIDTH-1:0] wire_d6_45;
	wire [WIDTH-1:0] wire_d6_46;
	wire [WIDTH-1:0] wire_d6_47;
	wire [WIDTH-1:0] wire_d6_48;
	wire [WIDTH-1:0] wire_d6_49;
	wire [WIDTH-1:0] wire_d6_50;
	wire [WIDTH-1:0] wire_d6_51;
	wire [WIDTH-1:0] wire_d6_52;
	wire [WIDTH-1:0] wire_d6_53;
	wire [WIDTH-1:0] wire_d6_54;
	wire [WIDTH-1:0] wire_d6_55;
	wire [WIDTH-1:0] wire_d6_56;
	wire [WIDTH-1:0] wire_d6_57;
	wire [WIDTH-1:0] wire_d6_58;
	wire [WIDTH-1:0] wire_d6_59;
	wire [WIDTH-1:0] wire_d6_60;
	wire [WIDTH-1:0] wire_d6_61;
	wire [WIDTH-1:0] wire_d6_62;
	wire [WIDTH-1:0] wire_d6_63;
	wire [WIDTH-1:0] wire_d6_64;
	wire [WIDTH-1:0] wire_d6_65;
	wire [WIDTH-1:0] wire_d6_66;
	wire [WIDTH-1:0] wire_d6_67;
	wire [WIDTH-1:0] wire_d6_68;
	wire [WIDTH-1:0] wire_d6_69;
	wire [WIDTH-1:0] wire_d6_70;
	wire [WIDTH-1:0] wire_d6_71;
	wire [WIDTH-1:0] wire_d6_72;
	wire [WIDTH-1:0] wire_d6_73;
	wire [WIDTH-1:0] wire_d6_74;
	wire [WIDTH-1:0] wire_d6_75;
	wire [WIDTH-1:0] wire_d6_76;
	wire [WIDTH-1:0] wire_d6_77;
	wire [WIDTH-1:0] wire_d6_78;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d7_29;
	wire [WIDTH-1:0] wire_d7_30;
	wire [WIDTH-1:0] wire_d7_31;
	wire [WIDTH-1:0] wire_d7_32;
	wire [WIDTH-1:0] wire_d7_33;
	wire [WIDTH-1:0] wire_d7_34;
	wire [WIDTH-1:0] wire_d7_35;
	wire [WIDTH-1:0] wire_d7_36;
	wire [WIDTH-1:0] wire_d7_37;
	wire [WIDTH-1:0] wire_d7_38;
	wire [WIDTH-1:0] wire_d7_39;
	wire [WIDTH-1:0] wire_d7_40;
	wire [WIDTH-1:0] wire_d7_41;
	wire [WIDTH-1:0] wire_d7_42;
	wire [WIDTH-1:0] wire_d7_43;
	wire [WIDTH-1:0] wire_d7_44;
	wire [WIDTH-1:0] wire_d7_45;
	wire [WIDTH-1:0] wire_d7_46;
	wire [WIDTH-1:0] wire_d7_47;
	wire [WIDTH-1:0] wire_d7_48;
	wire [WIDTH-1:0] wire_d7_49;
	wire [WIDTH-1:0] wire_d7_50;
	wire [WIDTH-1:0] wire_d7_51;
	wire [WIDTH-1:0] wire_d7_52;
	wire [WIDTH-1:0] wire_d7_53;
	wire [WIDTH-1:0] wire_d7_54;
	wire [WIDTH-1:0] wire_d7_55;
	wire [WIDTH-1:0] wire_d7_56;
	wire [WIDTH-1:0] wire_d7_57;
	wire [WIDTH-1:0] wire_d7_58;
	wire [WIDTH-1:0] wire_d7_59;
	wire [WIDTH-1:0] wire_d7_60;
	wire [WIDTH-1:0] wire_d7_61;
	wire [WIDTH-1:0] wire_d7_62;
	wire [WIDTH-1:0] wire_d7_63;
	wire [WIDTH-1:0] wire_d7_64;
	wire [WIDTH-1:0] wire_d7_65;
	wire [WIDTH-1:0] wire_d7_66;
	wire [WIDTH-1:0] wire_d7_67;
	wire [WIDTH-1:0] wire_d7_68;
	wire [WIDTH-1:0] wire_d7_69;
	wire [WIDTH-1:0] wire_d7_70;
	wire [WIDTH-1:0] wire_d7_71;
	wire [WIDTH-1:0] wire_d7_72;
	wire [WIDTH-1:0] wire_d7_73;
	wire [WIDTH-1:0] wire_d7_74;
	wire [WIDTH-1:0] wire_d7_75;
	wire [WIDTH-1:0] wire_d7_76;
	wire [WIDTH-1:0] wire_d7_77;
	wire [WIDTH-1:0] wire_d7_78;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d8_29;
	wire [WIDTH-1:0] wire_d8_30;
	wire [WIDTH-1:0] wire_d8_31;
	wire [WIDTH-1:0] wire_d8_32;
	wire [WIDTH-1:0] wire_d8_33;
	wire [WIDTH-1:0] wire_d8_34;
	wire [WIDTH-1:0] wire_d8_35;
	wire [WIDTH-1:0] wire_d8_36;
	wire [WIDTH-1:0] wire_d8_37;
	wire [WIDTH-1:0] wire_d8_38;
	wire [WIDTH-1:0] wire_d8_39;
	wire [WIDTH-1:0] wire_d8_40;
	wire [WIDTH-1:0] wire_d8_41;
	wire [WIDTH-1:0] wire_d8_42;
	wire [WIDTH-1:0] wire_d8_43;
	wire [WIDTH-1:0] wire_d8_44;
	wire [WIDTH-1:0] wire_d8_45;
	wire [WIDTH-1:0] wire_d8_46;
	wire [WIDTH-1:0] wire_d8_47;
	wire [WIDTH-1:0] wire_d8_48;
	wire [WIDTH-1:0] wire_d8_49;
	wire [WIDTH-1:0] wire_d8_50;
	wire [WIDTH-1:0] wire_d8_51;
	wire [WIDTH-1:0] wire_d8_52;
	wire [WIDTH-1:0] wire_d8_53;
	wire [WIDTH-1:0] wire_d8_54;
	wire [WIDTH-1:0] wire_d8_55;
	wire [WIDTH-1:0] wire_d8_56;
	wire [WIDTH-1:0] wire_d8_57;
	wire [WIDTH-1:0] wire_d8_58;
	wire [WIDTH-1:0] wire_d8_59;
	wire [WIDTH-1:0] wire_d8_60;
	wire [WIDTH-1:0] wire_d8_61;
	wire [WIDTH-1:0] wire_d8_62;
	wire [WIDTH-1:0] wire_d8_63;
	wire [WIDTH-1:0] wire_d8_64;
	wire [WIDTH-1:0] wire_d8_65;
	wire [WIDTH-1:0] wire_d8_66;
	wire [WIDTH-1:0] wire_d8_67;
	wire [WIDTH-1:0] wire_d8_68;
	wire [WIDTH-1:0] wire_d8_69;
	wire [WIDTH-1:0] wire_d8_70;
	wire [WIDTH-1:0] wire_d8_71;
	wire [WIDTH-1:0] wire_d8_72;
	wire [WIDTH-1:0] wire_d8_73;
	wire [WIDTH-1:0] wire_d8_74;
	wire [WIDTH-1:0] wire_d8_75;
	wire [WIDTH-1:0] wire_d8_76;
	wire [WIDTH-1:0] wire_d8_77;
	wire [WIDTH-1:0] wire_d8_78;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d9_29;
	wire [WIDTH-1:0] wire_d9_30;
	wire [WIDTH-1:0] wire_d9_31;
	wire [WIDTH-1:0] wire_d9_32;
	wire [WIDTH-1:0] wire_d9_33;
	wire [WIDTH-1:0] wire_d9_34;
	wire [WIDTH-1:0] wire_d9_35;
	wire [WIDTH-1:0] wire_d9_36;
	wire [WIDTH-1:0] wire_d9_37;
	wire [WIDTH-1:0] wire_d9_38;
	wire [WIDTH-1:0] wire_d9_39;
	wire [WIDTH-1:0] wire_d9_40;
	wire [WIDTH-1:0] wire_d9_41;
	wire [WIDTH-1:0] wire_d9_42;
	wire [WIDTH-1:0] wire_d9_43;
	wire [WIDTH-1:0] wire_d9_44;
	wire [WIDTH-1:0] wire_d9_45;
	wire [WIDTH-1:0] wire_d9_46;
	wire [WIDTH-1:0] wire_d9_47;
	wire [WIDTH-1:0] wire_d9_48;
	wire [WIDTH-1:0] wire_d9_49;
	wire [WIDTH-1:0] wire_d9_50;
	wire [WIDTH-1:0] wire_d9_51;
	wire [WIDTH-1:0] wire_d9_52;
	wire [WIDTH-1:0] wire_d9_53;
	wire [WIDTH-1:0] wire_d9_54;
	wire [WIDTH-1:0] wire_d9_55;
	wire [WIDTH-1:0] wire_d9_56;
	wire [WIDTH-1:0] wire_d9_57;
	wire [WIDTH-1:0] wire_d9_58;
	wire [WIDTH-1:0] wire_d9_59;
	wire [WIDTH-1:0] wire_d9_60;
	wire [WIDTH-1:0] wire_d9_61;
	wire [WIDTH-1:0] wire_d9_62;
	wire [WIDTH-1:0] wire_d9_63;
	wire [WIDTH-1:0] wire_d9_64;
	wire [WIDTH-1:0] wire_d9_65;
	wire [WIDTH-1:0] wire_d9_66;
	wire [WIDTH-1:0] wire_d9_67;
	wire [WIDTH-1:0] wire_d9_68;
	wire [WIDTH-1:0] wire_d9_69;
	wire [WIDTH-1:0] wire_d9_70;
	wire [WIDTH-1:0] wire_d9_71;
	wire [WIDTH-1:0] wire_d9_72;
	wire [WIDTH-1:0] wire_d9_73;
	wire [WIDTH-1:0] wire_d9_74;
	wire [WIDTH-1:0] wire_d9_75;
	wire [WIDTH-1:0] wire_d9_76;
	wire [WIDTH-1:0] wire_d9_77;
	wire [WIDTH-1:0] wire_d9_78;
	wire [WIDTH-1:0] wire_d10_0;
	wire [WIDTH-1:0] wire_d10_1;
	wire [WIDTH-1:0] wire_d10_2;
	wire [WIDTH-1:0] wire_d10_3;
	wire [WIDTH-1:0] wire_d10_4;
	wire [WIDTH-1:0] wire_d10_5;
	wire [WIDTH-1:0] wire_d10_6;
	wire [WIDTH-1:0] wire_d10_7;
	wire [WIDTH-1:0] wire_d10_8;
	wire [WIDTH-1:0] wire_d10_9;
	wire [WIDTH-1:0] wire_d10_10;
	wire [WIDTH-1:0] wire_d10_11;
	wire [WIDTH-1:0] wire_d10_12;
	wire [WIDTH-1:0] wire_d10_13;
	wire [WIDTH-1:0] wire_d10_14;
	wire [WIDTH-1:0] wire_d10_15;
	wire [WIDTH-1:0] wire_d10_16;
	wire [WIDTH-1:0] wire_d10_17;
	wire [WIDTH-1:0] wire_d10_18;
	wire [WIDTH-1:0] wire_d10_19;
	wire [WIDTH-1:0] wire_d10_20;
	wire [WIDTH-1:0] wire_d10_21;
	wire [WIDTH-1:0] wire_d10_22;
	wire [WIDTH-1:0] wire_d10_23;
	wire [WIDTH-1:0] wire_d10_24;
	wire [WIDTH-1:0] wire_d10_25;
	wire [WIDTH-1:0] wire_d10_26;
	wire [WIDTH-1:0] wire_d10_27;
	wire [WIDTH-1:0] wire_d10_28;
	wire [WIDTH-1:0] wire_d10_29;
	wire [WIDTH-1:0] wire_d10_30;
	wire [WIDTH-1:0] wire_d10_31;
	wire [WIDTH-1:0] wire_d10_32;
	wire [WIDTH-1:0] wire_d10_33;
	wire [WIDTH-1:0] wire_d10_34;
	wire [WIDTH-1:0] wire_d10_35;
	wire [WIDTH-1:0] wire_d10_36;
	wire [WIDTH-1:0] wire_d10_37;
	wire [WIDTH-1:0] wire_d10_38;
	wire [WIDTH-1:0] wire_d10_39;
	wire [WIDTH-1:0] wire_d10_40;
	wire [WIDTH-1:0] wire_d10_41;
	wire [WIDTH-1:0] wire_d10_42;
	wire [WIDTH-1:0] wire_d10_43;
	wire [WIDTH-1:0] wire_d10_44;
	wire [WIDTH-1:0] wire_d10_45;
	wire [WIDTH-1:0] wire_d10_46;
	wire [WIDTH-1:0] wire_d10_47;
	wire [WIDTH-1:0] wire_d10_48;
	wire [WIDTH-1:0] wire_d10_49;
	wire [WIDTH-1:0] wire_d10_50;
	wire [WIDTH-1:0] wire_d10_51;
	wire [WIDTH-1:0] wire_d10_52;
	wire [WIDTH-1:0] wire_d10_53;
	wire [WIDTH-1:0] wire_d10_54;
	wire [WIDTH-1:0] wire_d10_55;
	wire [WIDTH-1:0] wire_d10_56;
	wire [WIDTH-1:0] wire_d10_57;
	wire [WIDTH-1:0] wire_d10_58;
	wire [WIDTH-1:0] wire_d10_59;
	wire [WIDTH-1:0] wire_d10_60;
	wire [WIDTH-1:0] wire_d10_61;
	wire [WIDTH-1:0] wire_d10_62;
	wire [WIDTH-1:0] wire_d10_63;
	wire [WIDTH-1:0] wire_d10_64;
	wire [WIDTH-1:0] wire_d10_65;
	wire [WIDTH-1:0] wire_d10_66;
	wire [WIDTH-1:0] wire_d10_67;
	wire [WIDTH-1:0] wire_d10_68;
	wire [WIDTH-1:0] wire_d10_69;
	wire [WIDTH-1:0] wire_d10_70;
	wire [WIDTH-1:0] wire_d10_71;
	wire [WIDTH-1:0] wire_d10_72;
	wire [WIDTH-1:0] wire_d10_73;
	wire [WIDTH-1:0] wire_d10_74;
	wire [WIDTH-1:0] wire_d10_75;
	wire [WIDTH-1:0] wire_d10_76;
	wire [WIDTH-1:0] wire_d10_77;
	wire [WIDTH-1:0] wire_d10_78;
	wire [WIDTH-1:0] wire_d11_0;
	wire [WIDTH-1:0] wire_d11_1;
	wire [WIDTH-1:0] wire_d11_2;
	wire [WIDTH-1:0] wire_d11_3;
	wire [WIDTH-1:0] wire_d11_4;
	wire [WIDTH-1:0] wire_d11_5;
	wire [WIDTH-1:0] wire_d11_6;
	wire [WIDTH-1:0] wire_d11_7;
	wire [WIDTH-1:0] wire_d11_8;
	wire [WIDTH-1:0] wire_d11_9;
	wire [WIDTH-1:0] wire_d11_10;
	wire [WIDTH-1:0] wire_d11_11;
	wire [WIDTH-1:0] wire_d11_12;
	wire [WIDTH-1:0] wire_d11_13;
	wire [WIDTH-1:0] wire_d11_14;
	wire [WIDTH-1:0] wire_d11_15;
	wire [WIDTH-1:0] wire_d11_16;
	wire [WIDTH-1:0] wire_d11_17;
	wire [WIDTH-1:0] wire_d11_18;
	wire [WIDTH-1:0] wire_d11_19;
	wire [WIDTH-1:0] wire_d11_20;
	wire [WIDTH-1:0] wire_d11_21;
	wire [WIDTH-1:0] wire_d11_22;
	wire [WIDTH-1:0] wire_d11_23;
	wire [WIDTH-1:0] wire_d11_24;
	wire [WIDTH-1:0] wire_d11_25;
	wire [WIDTH-1:0] wire_d11_26;
	wire [WIDTH-1:0] wire_d11_27;
	wire [WIDTH-1:0] wire_d11_28;
	wire [WIDTH-1:0] wire_d11_29;
	wire [WIDTH-1:0] wire_d11_30;
	wire [WIDTH-1:0] wire_d11_31;
	wire [WIDTH-1:0] wire_d11_32;
	wire [WIDTH-1:0] wire_d11_33;
	wire [WIDTH-1:0] wire_d11_34;
	wire [WIDTH-1:0] wire_d11_35;
	wire [WIDTH-1:0] wire_d11_36;
	wire [WIDTH-1:0] wire_d11_37;
	wire [WIDTH-1:0] wire_d11_38;
	wire [WIDTH-1:0] wire_d11_39;
	wire [WIDTH-1:0] wire_d11_40;
	wire [WIDTH-1:0] wire_d11_41;
	wire [WIDTH-1:0] wire_d11_42;
	wire [WIDTH-1:0] wire_d11_43;
	wire [WIDTH-1:0] wire_d11_44;
	wire [WIDTH-1:0] wire_d11_45;
	wire [WIDTH-1:0] wire_d11_46;
	wire [WIDTH-1:0] wire_d11_47;
	wire [WIDTH-1:0] wire_d11_48;
	wire [WIDTH-1:0] wire_d11_49;
	wire [WIDTH-1:0] wire_d11_50;
	wire [WIDTH-1:0] wire_d11_51;
	wire [WIDTH-1:0] wire_d11_52;
	wire [WIDTH-1:0] wire_d11_53;
	wire [WIDTH-1:0] wire_d11_54;
	wire [WIDTH-1:0] wire_d11_55;
	wire [WIDTH-1:0] wire_d11_56;
	wire [WIDTH-1:0] wire_d11_57;
	wire [WIDTH-1:0] wire_d11_58;
	wire [WIDTH-1:0] wire_d11_59;
	wire [WIDTH-1:0] wire_d11_60;
	wire [WIDTH-1:0] wire_d11_61;
	wire [WIDTH-1:0] wire_d11_62;
	wire [WIDTH-1:0] wire_d11_63;
	wire [WIDTH-1:0] wire_d11_64;
	wire [WIDTH-1:0] wire_d11_65;
	wire [WIDTH-1:0] wire_d11_66;
	wire [WIDTH-1:0] wire_d11_67;
	wire [WIDTH-1:0] wire_d11_68;
	wire [WIDTH-1:0] wire_d11_69;
	wire [WIDTH-1:0] wire_d11_70;
	wire [WIDTH-1:0] wire_d11_71;
	wire [WIDTH-1:0] wire_d11_72;
	wire [WIDTH-1:0] wire_d11_73;
	wire [WIDTH-1:0] wire_d11_74;
	wire [WIDTH-1:0] wire_d11_75;
	wire [WIDTH-1:0] wire_d11_76;
	wire [WIDTH-1:0] wire_d11_77;
	wire [WIDTH-1:0] wire_d11_78;
	wire [WIDTH-1:0] wire_d12_0;
	wire [WIDTH-1:0] wire_d12_1;
	wire [WIDTH-1:0] wire_d12_2;
	wire [WIDTH-1:0] wire_d12_3;
	wire [WIDTH-1:0] wire_d12_4;
	wire [WIDTH-1:0] wire_d12_5;
	wire [WIDTH-1:0] wire_d12_6;
	wire [WIDTH-1:0] wire_d12_7;
	wire [WIDTH-1:0] wire_d12_8;
	wire [WIDTH-1:0] wire_d12_9;
	wire [WIDTH-1:0] wire_d12_10;
	wire [WIDTH-1:0] wire_d12_11;
	wire [WIDTH-1:0] wire_d12_12;
	wire [WIDTH-1:0] wire_d12_13;
	wire [WIDTH-1:0] wire_d12_14;
	wire [WIDTH-1:0] wire_d12_15;
	wire [WIDTH-1:0] wire_d12_16;
	wire [WIDTH-1:0] wire_d12_17;
	wire [WIDTH-1:0] wire_d12_18;
	wire [WIDTH-1:0] wire_d12_19;
	wire [WIDTH-1:0] wire_d12_20;
	wire [WIDTH-1:0] wire_d12_21;
	wire [WIDTH-1:0] wire_d12_22;
	wire [WIDTH-1:0] wire_d12_23;
	wire [WIDTH-1:0] wire_d12_24;
	wire [WIDTH-1:0] wire_d12_25;
	wire [WIDTH-1:0] wire_d12_26;
	wire [WIDTH-1:0] wire_d12_27;
	wire [WIDTH-1:0] wire_d12_28;
	wire [WIDTH-1:0] wire_d12_29;
	wire [WIDTH-1:0] wire_d12_30;
	wire [WIDTH-1:0] wire_d12_31;
	wire [WIDTH-1:0] wire_d12_32;
	wire [WIDTH-1:0] wire_d12_33;
	wire [WIDTH-1:0] wire_d12_34;
	wire [WIDTH-1:0] wire_d12_35;
	wire [WIDTH-1:0] wire_d12_36;
	wire [WIDTH-1:0] wire_d12_37;
	wire [WIDTH-1:0] wire_d12_38;
	wire [WIDTH-1:0] wire_d12_39;
	wire [WIDTH-1:0] wire_d12_40;
	wire [WIDTH-1:0] wire_d12_41;
	wire [WIDTH-1:0] wire_d12_42;
	wire [WIDTH-1:0] wire_d12_43;
	wire [WIDTH-1:0] wire_d12_44;
	wire [WIDTH-1:0] wire_d12_45;
	wire [WIDTH-1:0] wire_d12_46;
	wire [WIDTH-1:0] wire_d12_47;
	wire [WIDTH-1:0] wire_d12_48;
	wire [WIDTH-1:0] wire_d12_49;
	wire [WIDTH-1:0] wire_d12_50;
	wire [WIDTH-1:0] wire_d12_51;
	wire [WIDTH-1:0] wire_d12_52;
	wire [WIDTH-1:0] wire_d12_53;
	wire [WIDTH-1:0] wire_d12_54;
	wire [WIDTH-1:0] wire_d12_55;
	wire [WIDTH-1:0] wire_d12_56;
	wire [WIDTH-1:0] wire_d12_57;
	wire [WIDTH-1:0] wire_d12_58;
	wire [WIDTH-1:0] wire_d12_59;
	wire [WIDTH-1:0] wire_d12_60;
	wire [WIDTH-1:0] wire_d12_61;
	wire [WIDTH-1:0] wire_d12_62;
	wire [WIDTH-1:0] wire_d12_63;
	wire [WIDTH-1:0] wire_d12_64;
	wire [WIDTH-1:0] wire_d12_65;
	wire [WIDTH-1:0] wire_d12_66;
	wire [WIDTH-1:0] wire_d12_67;
	wire [WIDTH-1:0] wire_d12_68;
	wire [WIDTH-1:0] wire_d12_69;
	wire [WIDTH-1:0] wire_d12_70;
	wire [WIDTH-1:0] wire_d12_71;
	wire [WIDTH-1:0] wire_d12_72;
	wire [WIDTH-1:0] wire_d12_73;
	wire [WIDTH-1:0] wire_d12_74;
	wire [WIDTH-1:0] wire_d12_75;
	wire [WIDTH-1:0] wire_d12_76;
	wire [WIDTH-1:0] wire_d12_77;
	wire [WIDTH-1:0] wire_d12_78;
	wire [WIDTH-1:0] wire_d13_0;
	wire [WIDTH-1:0] wire_d13_1;
	wire [WIDTH-1:0] wire_d13_2;
	wire [WIDTH-1:0] wire_d13_3;
	wire [WIDTH-1:0] wire_d13_4;
	wire [WIDTH-1:0] wire_d13_5;
	wire [WIDTH-1:0] wire_d13_6;
	wire [WIDTH-1:0] wire_d13_7;
	wire [WIDTH-1:0] wire_d13_8;
	wire [WIDTH-1:0] wire_d13_9;
	wire [WIDTH-1:0] wire_d13_10;
	wire [WIDTH-1:0] wire_d13_11;
	wire [WIDTH-1:0] wire_d13_12;
	wire [WIDTH-1:0] wire_d13_13;
	wire [WIDTH-1:0] wire_d13_14;
	wire [WIDTH-1:0] wire_d13_15;
	wire [WIDTH-1:0] wire_d13_16;
	wire [WIDTH-1:0] wire_d13_17;
	wire [WIDTH-1:0] wire_d13_18;
	wire [WIDTH-1:0] wire_d13_19;
	wire [WIDTH-1:0] wire_d13_20;
	wire [WIDTH-1:0] wire_d13_21;
	wire [WIDTH-1:0] wire_d13_22;
	wire [WIDTH-1:0] wire_d13_23;
	wire [WIDTH-1:0] wire_d13_24;
	wire [WIDTH-1:0] wire_d13_25;
	wire [WIDTH-1:0] wire_d13_26;
	wire [WIDTH-1:0] wire_d13_27;
	wire [WIDTH-1:0] wire_d13_28;
	wire [WIDTH-1:0] wire_d13_29;
	wire [WIDTH-1:0] wire_d13_30;
	wire [WIDTH-1:0] wire_d13_31;
	wire [WIDTH-1:0] wire_d13_32;
	wire [WIDTH-1:0] wire_d13_33;
	wire [WIDTH-1:0] wire_d13_34;
	wire [WIDTH-1:0] wire_d13_35;
	wire [WIDTH-1:0] wire_d13_36;
	wire [WIDTH-1:0] wire_d13_37;
	wire [WIDTH-1:0] wire_d13_38;
	wire [WIDTH-1:0] wire_d13_39;
	wire [WIDTH-1:0] wire_d13_40;
	wire [WIDTH-1:0] wire_d13_41;
	wire [WIDTH-1:0] wire_d13_42;
	wire [WIDTH-1:0] wire_d13_43;
	wire [WIDTH-1:0] wire_d13_44;
	wire [WIDTH-1:0] wire_d13_45;
	wire [WIDTH-1:0] wire_d13_46;
	wire [WIDTH-1:0] wire_d13_47;
	wire [WIDTH-1:0] wire_d13_48;
	wire [WIDTH-1:0] wire_d13_49;
	wire [WIDTH-1:0] wire_d13_50;
	wire [WIDTH-1:0] wire_d13_51;
	wire [WIDTH-1:0] wire_d13_52;
	wire [WIDTH-1:0] wire_d13_53;
	wire [WIDTH-1:0] wire_d13_54;
	wire [WIDTH-1:0] wire_d13_55;
	wire [WIDTH-1:0] wire_d13_56;
	wire [WIDTH-1:0] wire_d13_57;
	wire [WIDTH-1:0] wire_d13_58;
	wire [WIDTH-1:0] wire_d13_59;
	wire [WIDTH-1:0] wire_d13_60;
	wire [WIDTH-1:0] wire_d13_61;
	wire [WIDTH-1:0] wire_d13_62;
	wire [WIDTH-1:0] wire_d13_63;
	wire [WIDTH-1:0] wire_d13_64;
	wire [WIDTH-1:0] wire_d13_65;
	wire [WIDTH-1:0] wire_d13_66;
	wire [WIDTH-1:0] wire_d13_67;
	wire [WIDTH-1:0] wire_d13_68;
	wire [WIDTH-1:0] wire_d13_69;
	wire [WIDTH-1:0] wire_d13_70;
	wire [WIDTH-1:0] wire_d13_71;
	wire [WIDTH-1:0] wire_d13_72;
	wire [WIDTH-1:0] wire_d13_73;
	wire [WIDTH-1:0] wire_d13_74;
	wire [WIDTH-1:0] wire_d13_75;
	wire [WIDTH-1:0] wire_d13_76;
	wire [WIDTH-1:0] wire_d13_77;
	wire [WIDTH-1:0] wire_d13_78;
	wire [WIDTH-1:0] wire_d14_0;
	wire [WIDTH-1:0] wire_d14_1;
	wire [WIDTH-1:0] wire_d14_2;
	wire [WIDTH-1:0] wire_d14_3;
	wire [WIDTH-1:0] wire_d14_4;
	wire [WIDTH-1:0] wire_d14_5;
	wire [WIDTH-1:0] wire_d14_6;
	wire [WIDTH-1:0] wire_d14_7;
	wire [WIDTH-1:0] wire_d14_8;
	wire [WIDTH-1:0] wire_d14_9;
	wire [WIDTH-1:0] wire_d14_10;
	wire [WIDTH-1:0] wire_d14_11;
	wire [WIDTH-1:0] wire_d14_12;
	wire [WIDTH-1:0] wire_d14_13;
	wire [WIDTH-1:0] wire_d14_14;
	wire [WIDTH-1:0] wire_d14_15;
	wire [WIDTH-1:0] wire_d14_16;
	wire [WIDTH-1:0] wire_d14_17;
	wire [WIDTH-1:0] wire_d14_18;
	wire [WIDTH-1:0] wire_d14_19;
	wire [WIDTH-1:0] wire_d14_20;
	wire [WIDTH-1:0] wire_d14_21;
	wire [WIDTH-1:0] wire_d14_22;
	wire [WIDTH-1:0] wire_d14_23;
	wire [WIDTH-1:0] wire_d14_24;
	wire [WIDTH-1:0] wire_d14_25;
	wire [WIDTH-1:0] wire_d14_26;
	wire [WIDTH-1:0] wire_d14_27;
	wire [WIDTH-1:0] wire_d14_28;
	wire [WIDTH-1:0] wire_d14_29;
	wire [WIDTH-1:0] wire_d14_30;
	wire [WIDTH-1:0] wire_d14_31;
	wire [WIDTH-1:0] wire_d14_32;
	wire [WIDTH-1:0] wire_d14_33;
	wire [WIDTH-1:0] wire_d14_34;
	wire [WIDTH-1:0] wire_d14_35;
	wire [WIDTH-1:0] wire_d14_36;
	wire [WIDTH-1:0] wire_d14_37;
	wire [WIDTH-1:0] wire_d14_38;
	wire [WIDTH-1:0] wire_d14_39;
	wire [WIDTH-1:0] wire_d14_40;
	wire [WIDTH-1:0] wire_d14_41;
	wire [WIDTH-1:0] wire_d14_42;
	wire [WIDTH-1:0] wire_d14_43;
	wire [WIDTH-1:0] wire_d14_44;
	wire [WIDTH-1:0] wire_d14_45;
	wire [WIDTH-1:0] wire_d14_46;
	wire [WIDTH-1:0] wire_d14_47;
	wire [WIDTH-1:0] wire_d14_48;
	wire [WIDTH-1:0] wire_d14_49;
	wire [WIDTH-1:0] wire_d14_50;
	wire [WIDTH-1:0] wire_d14_51;
	wire [WIDTH-1:0] wire_d14_52;
	wire [WIDTH-1:0] wire_d14_53;
	wire [WIDTH-1:0] wire_d14_54;
	wire [WIDTH-1:0] wire_d14_55;
	wire [WIDTH-1:0] wire_d14_56;
	wire [WIDTH-1:0] wire_d14_57;
	wire [WIDTH-1:0] wire_d14_58;
	wire [WIDTH-1:0] wire_d14_59;
	wire [WIDTH-1:0] wire_d14_60;
	wire [WIDTH-1:0] wire_d14_61;
	wire [WIDTH-1:0] wire_d14_62;
	wire [WIDTH-1:0] wire_d14_63;
	wire [WIDTH-1:0] wire_d14_64;
	wire [WIDTH-1:0] wire_d14_65;
	wire [WIDTH-1:0] wire_d14_66;
	wire [WIDTH-1:0] wire_d14_67;
	wire [WIDTH-1:0] wire_d14_68;
	wire [WIDTH-1:0] wire_d14_69;
	wire [WIDTH-1:0] wire_d14_70;
	wire [WIDTH-1:0] wire_d14_71;
	wire [WIDTH-1:0] wire_d14_72;
	wire [WIDTH-1:0] wire_d14_73;
	wire [WIDTH-1:0] wire_d14_74;
	wire [WIDTH-1:0] wire_d14_75;
	wire [WIDTH-1:0] wire_d14_76;
	wire [WIDTH-1:0] wire_d14_77;
	wire [WIDTH-1:0] wire_d14_78;
	wire [WIDTH-1:0] wire_d15_0;
	wire [WIDTH-1:0] wire_d15_1;
	wire [WIDTH-1:0] wire_d15_2;
	wire [WIDTH-1:0] wire_d15_3;
	wire [WIDTH-1:0] wire_d15_4;
	wire [WIDTH-1:0] wire_d15_5;
	wire [WIDTH-1:0] wire_d15_6;
	wire [WIDTH-1:0] wire_d15_7;
	wire [WIDTH-1:0] wire_d15_8;
	wire [WIDTH-1:0] wire_d15_9;
	wire [WIDTH-1:0] wire_d15_10;
	wire [WIDTH-1:0] wire_d15_11;
	wire [WIDTH-1:0] wire_d15_12;
	wire [WIDTH-1:0] wire_d15_13;
	wire [WIDTH-1:0] wire_d15_14;
	wire [WIDTH-1:0] wire_d15_15;
	wire [WIDTH-1:0] wire_d15_16;
	wire [WIDTH-1:0] wire_d15_17;
	wire [WIDTH-1:0] wire_d15_18;
	wire [WIDTH-1:0] wire_d15_19;
	wire [WIDTH-1:0] wire_d15_20;
	wire [WIDTH-1:0] wire_d15_21;
	wire [WIDTH-1:0] wire_d15_22;
	wire [WIDTH-1:0] wire_d15_23;
	wire [WIDTH-1:0] wire_d15_24;
	wire [WIDTH-1:0] wire_d15_25;
	wire [WIDTH-1:0] wire_d15_26;
	wire [WIDTH-1:0] wire_d15_27;
	wire [WIDTH-1:0] wire_d15_28;
	wire [WIDTH-1:0] wire_d15_29;
	wire [WIDTH-1:0] wire_d15_30;
	wire [WIDTH-1:0] wire_d15_31;
	wire [WIDTH-1:0] wire_d15_32;
	wire [WIDTH-1:0] wire_d15_33;
	wire [WIDTH-1:0] wire_d15_34;
	wire [WIDTH-1:0] wire_d15_35;
	wire [WIDTH-1:0] wire_d15_36;
	wire [WIDTH-1:0] wire_d15_37;
	wire [WIDTH-1:0] wire_d15_38;
	wire [WIDTH-1:0] wire_d15_39;
	wire [WIDTH-1:0] wire_d15_40;
	wire [WIDTH-1:0] wire_d15_41;
	wire [WIDTH-1:0] wire_d15_42;
	wire [WIDTH-1:0] wire_d15_43;
	wire [WIDTH-1:0] wire_d15_44;
	wire [WIDTH-1:0] wire_d15_45;
	wire [WIDTH-1:0] wire_d15_46;
	wire [WIDTH-1:0] wire_d15_47;
	wire [WIDTH-1:0] wire_d15_48;
	wire [WIDTH-1:0] wire_d15_49;
	wire [WIDTH-1:0] wire_d15_50;
	wire [WIDTH-1:0] wire_d15_51;
	wire [WIDTH-1:0] wire_d15_52;
	wire [WIDTH-1:0] wire_d15_53;
	wire [WIDTH-1:0] wire_d15_54;
	wire [WIDTH-1:0] wire_d15_55;
	wire [WIDTH-1:0] wire_d15_56;
	wire [WIDTH-1:0] wire_d15_57;
	wire [WIDTH-1:0] wire_d15_58;
	wire [WIDTH-1:0] wire_d15_59;
	wire [WIDTH-1:0] wire_d15_60;
	wire [WIDTH-1:0] wire_d15_61;
	wire [WIDTH-1:0] wire_d15_62;
	wire [WIDTH-1:0] wire_d15_63;
	wire [WIDTH-1:0] wire_d15_64;
	wire [WIDTH-1:0] wire_d15_65;
	wire [WIDTH-1:0] wire_d15_66;
	wire [WIDTH-1:0] wire_d15_67;
	wire [WIDTH-1:0] wire_d15_68;
	wire [WIDTH-1:0] wire_d15_69;
	wire [WIDTH-1:0] wire_d15_70;
	wire [WIDTH-1:0] wire_d15_71;
	wire [WIDTH-1:0] wire_d15_72;
	wire [WIDTH-1:0] wire_d15_73;
	wire [WIDTH-1:0] wire_d15_74;
	wire [WIDTH-1:0] wire_d15_75;
	wire [WIDTH-1:0] wire_d15_76;
	wire [WIDTH-1:0] wire_d15_77;
	wire [WIDTH-1:0] wire_d15_78;
	wire [WIDTH-1:0] wire_d16_0;
	wire [WIDTH-1:0] wire_d16_1;
	wire [WIDTH-1:0] wire_d16_2;
	wire [WIDTH-1:0] wire_d16_3;
	wire [WIDTH-1:0] wire_d16_4;
	wire [WIDTH-1:0] wire_d16_5;
	wire [WIDTH-1:0] wire_d16_6;
	wire [WIDTH-1:0] wire_d16_7;
	wire [WIDTH-1:0] wire_d16_8;
	wire [WIDTH-1:0] wire_d16_9;
	wire [WIDTH-1:0] wire_d16_10;
	wire [WIDTH-1:0] wire_d16_11;
	wire [WIDTH-1:0] wire_d16_12;
	wire [WIDTH-1:0] wire_d16_13;
	wire [WIDTH-1:0] wire_d16_14;
	wire [WIDTH-1:0] wire_d16_15;
	wire [WIDTH-1:0] wire_d16_16;
	wire [WIDTH-1:0] wire_d16_17;
	wire [WIDTH-1:0] wire_d16_18;
	wire [WIDTH-1:0] wire_d16_19;
	wire [WIDTH-1:0] wire_d16_20;
	wire [WIDTH-1:0] wire_d16_21;
	wire [WIDTH-1:0] wire_d16_22;
	wire [WIDTH-1:0] wire_d16_23;
	wire [WIDTH-1:0] wire_d16_24;
	wire [WIDTH-1:0] wire_d16_25;
	wire [WIDTH-1:0] wire_d16_26;
	wire [WIDTH-1:0] wire_d16_27;
	wire [WIDTH-1:0] wire_d16_28;
	wire [WIDTH-1:0] wire_d16_29;
	wire [WIDTH-1:0] wire_d16_30;
	wire [WIDTH-1:0] wire_d16_31;
	wire [WIDTH-1:0] wire_d16_32;
	wire [WIDTH-1:0] wire_d16_33;
	wire [WIDTH-1:0] wire_d16_34;
	wire [WIDTH-1:0] wire_d16_35;
	wire [WIDTH-1:0] wire_d16_36;
	wire [WIDTH-1:0] wire_d16_37;
	wire [WIDTH-1:0] wire_d16_38;
	wire [WIDTH-1:0] wire_d16_39;
	wire [WIDTH-1:0] wire_d16_40;
	wire [WIDTH-1:0] wire_d16_41;
	wire [WIDTH-1:0] wire_d16_42;
	wire [WIDTH-1:0] wire_d16_43;
	wire [WIDTH-1:0] wire_d16_44;
	wire [WIDTH-1:0] wire_d16_45;
	wire [WIDTH-1:0] wire_d16_46;
	wire [WIDTH-1:0] wire_d16_47;
	wire [WIDTH-1:0] wire_d16_48;
	wire [WIDTH-1:0] wire_d16_49;
	wire [WIDTH-1:0] wire_d16_50;
	wire [WIDTH-1:0] wire_d16_51;
	wire [WIDTH-1:0] wire_d16_52;
	wire [WIDTH-1:0] wire_d16_53;
	wire [WIDTH-1:0] wire_d16_54;
	wire [WIDTH-1:0] wire_d16_55;
	wire [WIDTH-1:0] wire_d16_56;
	wire [WIDTH-1:0] wire_d16_57;
	wire [WIDTH-1:0] wire_d16_58;
	wire [WIDTH-1:0] wire_d16_59;
	wire [WIDTH-1:0] wire_d16_60;
	wire [WIDTH-1:0] wire_d16_61;
	wire [WIDTH-1:0] wire_d16_62;
	wire [WIDTH-1:0] wire_d16_63;
	wire [WIDTH-1:0] wire_d16_64;
	wire [WIDTH-1:0] wire_d16_65;
	wire [WIDTH-1:0] wire_d16_66;
	wire [WIDTH-1:0] wire_d16_67;
	wire [WIDTH-1:0] wire_d16_68;
	wire [WIDTH-1:0] wire_d16_69;
	wire [WIDTH-1:0] wire_d16_70;
	wire [WIDTH-1:0] wire_d16_71;
	wire [WIDTH-1:0] wire_d16_72;
	wire [WIDTH-1:0] wire_d16_73;
	wire [WIDTH-1:0] wire_d16_74;
	wire [WIDTH-1:0] wire_d16_75;
	wire [WIDTH-1:0] wire_d16_76;
	wire [WIDTH-1:0] wire_d16_77;
	wire [WIDTH-1:0] wire_d16_78;
	wire [WIDTH-1:0] wire_d17_0;
	wire [WIDTH-1:0] wire_d17_1;
	wire [WIDTH-1:0] wire_d17_2;
	wire [WIDTH-1:0] wire_d17_3;
	wire [WIDTH-1:0] wire_d17_4;
	wire [WIDTH-1:0] wire_d17_5;
	wire [WIDTH-1:0] wire_d17_6;
	wire [WIDTH-1:0] wire_d17_7;
	wire [WIDTH-1:0] wire_d17_8;
	wire [WIDTH-1:0] wire_d17_9;
	wire [WIDTH-1:0] wire_d17_10;
	wire [WIDTH-1:0] wire_d17_11;
	wire [WIDTH-1:0] wire_d17_12;
	wire [WIDTH-1:0] wire_d17_13;
	wire [WIDTH-1:0] wire_d17_14;
	wire [WIDTH-1:0] wire_d17_15;
	wire [WIDTH-1:0] wire_d17_16;
	wire [WIDTH-1:0] wire_d17_17;
	wire [WIDTH-1:0] wire_d17_18;
	wire [WIDTH-1:0] wire_d17_19;
	wire [WIDTH-1:0] wire_d17_20;
	wire [WIDTH-1:0] wire_d17_21;
	wire [WIDTH-1:0] wire_d17_22;
	wire [WIDTH-1:0] wire_d17_23;
	wire [WIDTH-1:0] wire_d17_24;
	wire [WIDTH-1:0] wire_d17_25;
	wire [WIDTH-1:0] wire_d17_26;
	wire [WIDTH-1:0] wire_d17_27;
	wire [WIDTH-1:0] wire_d17_28;
	wire [WIDTH-1:0] wire_d17_29;
	wire [WIDTH-1:0] wire_d17_30;
	wire [WIDTH-1:0] wire_d17_31;
	wire [WIDTH-1:0] wire_d17_32;
	wire [WIDTH-1:0] wire_d17_33;
	wire [WIDTH-1:0] wire_d17_34;
	wire [WIDTH-1:0] wire_d17_35;
	wire [WIDTH-1:0] wire_d17_36;
	wire [WIDTH-1:0] wire_d17_37;
	wire [WIDTH-1:0] wire_d17_38;
	wire [WIDTH-1:0] wire_d17_39;
	wire [WIDTH-1:0] wire_d17_40;
	wire [WIDTH-1:0] wire_d17_41;
	wire [WIDTH-1:0] wire_d17_42;
	wire [WIDTH-1:0] wire_d17_43;
	wire [WIDTH-1:0] wire_d17_44;
	wire [WIDTH-1:0] wire_d17_45;
	wire [WIDTH-1:0] wire_d17_46;
	wire [WIDTH-1:0] wire_d17_47;
	wire [WIDTH-1:0] wire_d17_48;
	wire [WIDTH-1:0] wire_d17_49;
	wire [WIDTH-1:0] wire_d17_50;
	wire [WIDTH-1:0] wire_d17_51;
	wire [WIDTH-1:0] wire_d17_52;
	wire [WIDTH-1:0] wire_d17_53;
	wire [WIDTH-1:0] wire_d17_54;
	wire [WIDTH-1:0] wire_d17_55;
	wire [WIDTH-1:0] wire_d17_56;
	wire [WIDTH-1:0] wire_d17_57;
	wire [WIDTH-1:0] wire_d17_58;
	wire [WIDTH-1:0] wire_d17_59;
	wire [WIDTH-1:0] wire_d17_60;
	wire [WIDTH-1:0] wire_d17_61;
	wire [WIDTH-1:0] wire_d17_62;
	wire [WIDTH-1:0] wire_d17_63;
	wire [WIDTH-1:0] wire_d17_64;
	wire [WIDTH-1:0] wire_d17_65;
	wire [WIDTH-1:0] wire_d17_66;
	wire [WIDTH-1:0] wire_d17_67;
	wire [WIDTH-1:0] wire_d17_68;
	wire [WIDTH-1:0] wire_d17_69;
	wire [WIDTH-1:0] wire_d17_70;
	wire [WIDTH-1:0] wire_d17_71;
	wire [WIDTH-1:0] wire_d17_72;
	wire [WIDTH-1:0] wire_d17_73;
	wire [WIDTH-1:0] wire_d17_74;
	wire [WIDTH-1:0] wire_d17_75;
	wire [WIDTH-1:0] wire_d17_76;
	wire [WIDTH-1:0] wire_d17_77;
	wire [WIDTH-1:0] wire_d17_78;
	wire [WIDTH-1:0] wire_d18_0;
	wire [WIDTH-1:0] wire_d18_1;
	wire [WIDTH-1:0] wire_d18_2;
	wire [WIDTH-1:0] wire_d18_3;
	wire [WIDTH-1:0] wire_d18_4;
	wire [WIDTH-1:0] wire_d18_5;
	wire [WIDTH-1:0] wire_d18_6;
	wire [WIDTH-1:0] wire_d18_7;
	wire [WIDTH-1:0] wire_d18_8;
	wire [WIDTH-1:0] wire_d18_9;
	wire [WIDTH-1:0] wire_d18_10;
	wire [WIDTH-1:0] wire_d18_11;
	wire [WIDTH-1:0] wire_d18_12;
	wire [WIDTH-1:0] wire_d18_13;
	wire [WIDTH-1:0] wire_d18_14;
	wire [WIDTH-1:0] wire_d18_15;
	wire [WIDTH-1:0] wire_d18_16;
	wire [WIDTH-1:0] wire_d18_17;
	wire [WIDTH-1:0] wire_d18_18;
	wire [WIDTH-1:0] wire_d18_19;
	wire [WIDTH-1:0] wire_d18_20;
	wire [WIDTH-1:0] wire_d18_21;
	wire [WIDTH-1:0] wire_d18_22;
	wire [WIDTH-1:0] wire_d18_23;
	wire [WIDTH-1:0] wire_d18_24;
	wire [WIDTH-1:0] wire_d18_25;
	wire [WIDTH-1:0] wire_d18_26;
	wire [WIDTH-1:0] wire_d18_27;
	wire [WIDTH-1:0] wire_d18_28;
	wire [WIDTH-1:0] wire_d18_29;
	wire [WIDTH-1:0] wire_d18_30;
	wire [WIDTH-1:0] wire_d18_31;
	wire [WIDTH-1:0] wire_d18_32;
	wire [WIDTH-1:0] wire_d18_33;
	wire [WIDTH-1:0] wire_d18_34;
	wire [WIDTH-1:0] wire_d18_35;
	wire [WIDTH-1:0] wire_d18_36;
	wire [WIDTH-1:0] wire_d18_37;
	wire [WIDTH-1:0] wire_d18_38;
	wire [WIDTH-1:0] wire_d18_39;
	wire [WIDTH-1:0] wire_d18_40;
	wire [WIDTH-1:0] wire_d18_41;
	wire [WIDTH-1:0] wire_d18_42;
	wire [WIDTH-1:0] wire_d18_43;
	wire [WIDTH-1:0] wire_d18_44;
	wire [WIDTH-1:0] wire_d18_45;
	wire [WIDTH-1:0] wire_d18_46;
	wire [WIDTH-1:0] wire_d18_47;
	wire [WIDTH-1:0] wire_d18_48;
	wire [WIDTH-1:0] wire_d18_49;
	wire [WIDTH-1:0] wire_d18_50;
	wire [WIDTH-1:0] wire_d18_51;
	wire [WIDTH-1:0] wire_d18_52;
	wire [WIDTH-1:0] wire_d18_53;
	wire [WIDTH-1:0] wire_d18_54;
	wire [WIDTH-1:0] wire_d18_55;
	wire [WIDTH-1:0] wire_d18_56;
	wire [WIDTH-1:0] wire_d18_57;
	wire [WIDTH-1:0] wire_d18_58;
	wire [WIDTH-1:0] wire_d18_59;
	wire [WIDTH-1:0] wire_d18_60;
	wire [WIDTH-1:0] wire_d18_61;
	wire [WIDTH-1:0] wire_d18_62;
	wire [WIDTH-1:0] wire_d18_63;
	wire [WIDTH-1:0] wire_d18_64;
	wire [WIDTH-1:0] wire_d18_65;
	wire [WIDTH-1:0] wire_d18_66;
	wire [WIDTH-1:0] wire_d18_67;
	wire [WIDTH-1:0] wire_d18_68;
	wire [WIDTH-1:0] wire_d18_69;
	wire [WIDTH-1:0] wire_d18_70;
	wire [WIDTH-1:0] wire_d18_71;
	wire [WIDTH-1:0] wire_d18_72;
	wire [WIDTH-1:0] wire_d18_73;
	wire [WIDTH-1:0] wire_d18_74;
	wire [WIDTH-1:0] wire_d18_75;
	wire [WIDTH-1:0] wire_d18_76;
	wire [WIDTH-1:0] wire_d18_77;
	wire [WIDTH-1:0] wire_d18_78;
	wire [WIDTH-1:0] wire_d19_0;
	wire [WIDTH-1:0] wire_d19_1;
	wire [WIDTH-1:0] wire_d19_2;
	wire [WIDTH-1:0] wire_d19_3;
	wire [WIDTH-1:0] wire_d19_4;
	wire [WIDTH-1:0] wire_d19_5;
	wire [WIDTH-1:0] wire_d19_6;
	wire [WIDTH-1:0] wire_d19_7;
	wire [WIDTH-1:0] wire_d19_8;
	wire [WIDTH-1:0] wire_d19_9;
	wire [WIDTH-1:0] wire_d19_10;
	wire [WIDTH-1:0] wire_d19_11;
	wire [WIDTH-1:0] wire_d19_12;
	wire [WIDTH-1:0] wire_d19_13;
	wire [WIDTH-1:0] wire_d19_14;
	wire [WIDTH-1:0] wire_d19_15;
	wire [WIDTH-1:0] wire_d19_16;
	wire [WIDTH-1:0] wire_d19_17;
	wire [WIDTH-1:0] wire_d19_18;
	wire [WIDTH-1:0] wire_d19_19;
	wire [WIDTH-1:0] wire_d19_20;
	wire [WIDTH-1:0] wire_d19_21;
	wire [WIDTH-1:0] wire_d19_22;
	wire [WIDTH-1:0] wire_d19_23;
	wire [WIDTH-1:0] wire_d19_24;
	wire [WIDTH-1:0] wire_d19_25;
	wire [WIDTH-1:0] wire_d19_26;
	wire [WIDTH-1:0] wire_d19_27;
	wire [WIDTH-1:0] wire_d19_28;
	wire [WIDTH-1:0] wire_d19_29;
	wire [WIDTH-1:0] wire_d19_30;
	wire [WIDTH-1:0] wire_d19_31;
	wire [WIDTH-1:0] wire_d19_32;
	wire [WIDTH-1:0] wire_d19_33;
	wire [WIDTH-1:0] wire_d19_34;
	wire [WIDTH-1:0] wire_d19_35;
	wire [WIDTH-1:0] wire_d19_36;
	wire [WIDTH-1:0] wire_d19_37;
	wire [WIDTH-1:0] wire_d19_38;
	wire [WIDTH-1:0] wire_d19_39;
	wire [WIDTH-1:0] wire_d19_40;
	wire [WIDTH-1:0] wire_d19_41;
	wire [WIDTH-1:0] wire_d19_42;
	wire [WIDTH-1:0] wire_d19_43;
	wire [WIDTH-1:0] wire_d19_44;
	wire [WIDTH-1:0] wire_d19_45;
	wire [WIDTH-1:0] wire_d19_46;
	wire [WIDTH-1:0] wire_d19_47;
	wire [WIDTH-1:0] wire_d19_48;
	wire [WIDTH-1:0] wire_d19_49;
	wire [WIDTH-1:0] wire_d19_50;
	wire [WIDTH-1:0] wire_d19_51;
	wire [WIDTH-1:0] wire_d19_52;
	wire [WIDTH-1:0] wire_d19_53;
	wire [WIDTH-1:0] wire_d19_54;
	wire [WIDTH-1:0] wire_d19_55;
	wire [WIDTH-1:0] wire_d19_56;
	wire [WIDTH-1:0] wire_d19_57;
	wire [WIDTH-1:0] wire_d19_58;
	wire [WIDTH-1:0] wire_d19_59;
	wire [WIDTH-1:0] wire_d19_60;
	wire [WIDTH-1:0] wire_d19_61;
	wire [WIDTH-1:0] wire_d19_62;
	wire [WIDTH-1:0] wire_d19_63;
	wire [WIDTH-1:0] wire_d19_64;
	wire [WIDTH-1:0] wire_d19_65;
	wire [WIDTH-1:0] wire_d19_66;
	wire [WIDTH-1:0] wire_d19_67;
	wire [WIDTH-1:0] wire_d19_68;
	wire [WIDTH-1:0] wire_d19_69;
	wire [WIDTH-1:0] wire_d19_70;
	wire [WIDTH-1:0] wire_d19_71;
	wire [WIDTH-1:0] wire_d19_72;
	wire [WIDTH-1:0] wire_d19_73;
	wire [WIDTH-1:0] wire_d19_74;
	wire [WIDTH-1:0] wire_d19_75;
	wire [WIDTH-1:0] wire_d19_76;
	wire [WIDTH-1:0] wire_d19_77;
	wire [WIDTH-1:0] wire_d19_78;
	wire [WIDTH-1:0] wire_d20_0;
	wire [WIDTH-1:0] wire_d20_1;
	wire [WIDTH-1:0] wire_d20_2;
	wire [WIDTH-1:0] wire_d20_3;
	wire [WIDTH-1:0] wire_d20_4;
	wire [WIDTH-1:0] wire_d20_5;
	wire [WIDTH-1:0] wire_d20_6;
	wire [WIDTH-1:0] wire_d20_7;
	wire [WIDTH-1:0] wire_d20_8;
	wire [WIDTH-1:0] wire_d20_9;
	wire [WIDTH-1:0] wire_d20_10;
	wire [WIDTH-1:0] wire_d20_11;
	wire [WIDTH-1:0] wire_d20_12;
	wire [WIDTH-1:0] wire_d20_13;
	wire [WIDTH-1:0] wire_d20_14;
	wire [WIDTH-1:0] wire_d20_15;
	wire [WIDTH-1:0] wire_d20_16;
	wire [WIDTH-1:0] wire_d20_17;
	wire [WIDTH-1:0] wire_d20_18;
	wire [WIDTH-1:0] wire_d20_19;
	wire [WIDTH-1:0] wire_d20_20;
	wire [WIDTH-1:0] wire_d20_21;
	wire [WIDTH-1:0] wire_d20_22;
	wire [WIDTH-1:0] wire_d20_23;
	wire [WIDTH-1:0] wire_d20_24;
	wire [WIDTH-1:0] wire_d20_25;
	wire [WIDTH-1:0] wire_d20_26;
	wire [WIDTH-1:0] wire_d20_27;
	wire [WIDTH-1:0] wire_d20_28;
	wire [WIDTH-1:0] wire_d20_29;
	wire [WIDTH-1:0] wire_d20_30;
	wire [WIDTH-1:0] wire_d20_31;
	wire [WIDTH-1:0] wire_d20_32;
	wire [WIDTH-1:0] wire_d20_33;
	wire [WIDTH-1:0] wire_d20_34;
	wire [WIDTH-1:0] wire_d20_35;
	wire [WIDTH-1:0] wire_d20_36;
	wire [WIDTH-1:0] wire_d20_37;
	wire [WIDTH-1:0] wire_d20_38;
	wire [WIDTH-1:0] wire_d20_39;
	wire [WIDTH-1:0] wire_d20_40;
	wire [WIDTH-1:0] wire_d20_41;
	wire [WIDTH-1:0] wire_d20_42;
	wire [WIDTH-1:0] wire_d20_43;
	wire [WIDTH-1:0] wire_d20_44;
	wire [WIDTH-1:0] wire_d20_45;
	wire [WIDTH-1:0] wire_d20_46;
	wire [WIDTH-1:0] wire_d20_47;
	wire [WIDTH-1:0] wire_d20_48;
	wire [WIDTH-1:0] wire_d20_49;
	wire [WIDTH-1:0] wire_d20_50;
	wire [WIDTH-1:0] wire_d20_51;
	wire [WIDTH-1:0] wire_d20_52;
	wire [WIDTH-1:0] wire_d20_53;
	wire [WIDTH-1:0] wire_d20_54;
	wire [WIDTH-1:0] wire_d20_55;
	wire [WIDTH-1:0] wire_d20_56;
	wire [WIDTH-1:0] wire_d20_57;
	wire [WIDTH-1:0] wire_d20_58;
	wire [WIDTH-1:0] wire_d20_59;
	wire [WIDTH-1:0] wire_d20_60;
	wire [WIDTH-1:0] wire_d20_61;
	wire [WIDTH-1:0] wire_d20_62;
	wire [WIDTH-1:0] wire_d20_63;
	wire [WIDTH-1:0] wire_d20_64;
	wire [WIDTH-1:0] wire_d20_65;
	wire [WIDTH-1:0] wire_d20_66;
	wire [WIDTH-1:0] wire_d20_67;
	wire [WIDTH-1:0] wire_d20_68;
	wire [WIDTH-1:0] wire_d20_69;
	wire [WIDTH-1:0] wire_d20_70;
	wire [WIDTH-1:0] wire_d20_71;
	wire [WIDTH-1:0] wire_d20_72;
	wire [WIDTH-1:0] wire_d20_73;
	wire [WIDTH-1:0] wire_d20_74;
	wire [WIDTH-1:0] wire_d20_75;
	wire [WIDTH-1:0] wire_d20_76;
	wire [WIDTH-1:0] wire_d20_77;
	wire [WIDTH-1:0] wire_d20_78;
	wire [WIDTH-1:0] wire_d21_0;
	wire [WIDTH-1:0] wire_d21_1;
	wire [WIDTH-1:0] wire_d21_2;
	wire [WIDTH-1:0] wire_d21_3;
	wire [WIDTH-1:0] wire_d21_4;
	wire [WIDTH-1:0] wire_d21_5;
	wire [WIDTH-1:0] wire_d21_6;
	wire [WIDTH-1:0] wire_d21_7;
	wire [WIDTH-1:0] wire_d21_8;
	wire [WIDTH-1:0] wire_d21_9;
	wire [WIDTH-1:0] wire_d21_10;
	wire [WIDTH-1:0] wire_d21_11;
	wire [WIDTH-1:0] wire_d21_12;
	wire [WIDTH-1:0] wire_d21_13;
	wire [WIDTH-1:0] wire_d21_14;
	wire [WIDTH-1:0] wire_d21_15;
	wire [WIDTH-1:0] wire_d21_16;
	wire [WIDTH-1:0] wire_d21_17;
	wire [WIDTH-1:0] wire_d21_18;
	wire [WIDTH-1:0] wire_d21_19;
	wire [WIDTH-1:0] wire_d21_20;
	wire [WIDTH-1:0] wire_d21_21;
	wire [WIDTH-1:0] wire_d21_22;
	wire [WIDTH-1:0] wire_d21_23;
	wire [WIDTH-1:0] wire_d21_24;
	wire [WIDTH-1:0] wire_d21_25;
	wire [WIDTH-1:0] wire_d21_26;
	wire [WIDTH-1:0] wire_d21_27;
	wire [WIDTH-1:0] wire_d21_28;
	wire [WIDTH-1:0] wire_d21_29;
	wire [WIDTH-1:0] wire_d21_30;
	wire [WIDTH-1:0] wire_d21_31;
	wire [WIDTH-1:0] wire_d21_32;
	wire [WIDTH-1:0] wire_d21_33;
	wire [WIDTH-1:0] wire_d21_34;
	wire [WIDTH-1:0] wire_d21_35;
	wire [WIDTH-1:0] wire_d21_36;
	wire [WIDTH-1:0] wire_d21_37;
	wire [WIDTH-1:0] wire_d21_38;
	wire [WIDTH-1:0] wire_d21_39;
	wire [WIDTH-1:0] wire_d21_40;
	wire [WIDTH-1:0] wire_d21_41;
	wire [WIDTH-1:0] wire_d21_42;
	wire [WIDTH-1:0] wire_d21_43;
	wire [WIDTH-1:0] wire_d21_44;
	wire [WIDTH-1:0] wire_d21_45;
	wire [WIDTH-1:0] wire_d21_46;
	wire [WIDTH-1:0] wire_d21_47;
	wire [WIDTH-1:0] wire_d21_48;
	wire [WIDTH-1:0] wire_d21_49;
	wire [WIDTH-1:0] wire_d21_50;
	wire [WIDTH-1:0] wire_d21_51;
	wire [WIDTH-1:0] wire_d21_52;
	wire [WIDTH-1:0] wire_d21_53;
	wire [WIDTH-1:0] wire_d21_54;
	wire [WIDTH-1:0] wire_d21_55;
	wire [WIDTH-1:0] wire_d21_56;
	wire [WIDTH-1:0] wire_d21_57;
	wire [WIDTH-1:0] wire_d21_58;
	wire [WIDTH-1:0] wire_d21_59;
	wire [WIDTH-1:0] wire_d21_60;
	wire [WIDTH-1:0] wire_d21_61;
	wire [WIDTH-1:0] wire_d21_62;
	wire [WIDTH-1:0] wire_d21_63;
	wire [WIDTH-1:0] wire_d21_64;
	wire [WIDTH-1:0] wire_d21_65;
	wire [WIDTH-1:0] wire_d21_66;
	wire [WIDTH-1:0] wire_d21_67;
	wire [WIDTH-1:0] wire_d21_68;
	wire [WIDTH-1:0] wire_d21_69;
	wire [WIDTH-1:0] wire_d21_70;
	wire [WIDTH-1:0] wire_d21_71;
	wire [WIDTH-1:0] wire_d21_72;
	wire [WIDTH-1:0] wire_d21_73;
	wire [WIDTH-1:0] wire_d21_74;
	wire [WIDTH-1:0] wire_d21_75;
	wire [WIDTH-1:0] wire_d21_76;
	wire [WIDTH-1:0] wire_d21_77;
	wire [WIDTH-1:0] wire_d21_78;
	wire [WIDTH-1:0] wire_d22_0;
	wire [WIDTH-1:0] wire_d22_1;
	wire [WIDTH-1:0] wire_d22_2;
	wire [WIDTH-1:0] wire_d22_3;
	wire [WIDTH-1:0] wire_d22_4;
	wire [WIDTH-1:0] wire_d22_5;
	wire [WIDTH-1:0] wire_d22_6;
	wire [WIDTH-1:0] wire_d22_7;
	wire [WIDTH-1:0] wire_d22_8;
	wire [WIDTH-1:0] wire_d22_9;
	wire [WIDTH-1:0] wire_d22_10;
	wire [WIDTH-1:0] wire_d22_11;
	wire [WIDTH-1:0] wire_d22_12;
	wire [WIDTH-1:0] wire_d22_13;
	wire [WIDTH-1:0] wire_d22_14;
	wire [WIDTH-1:0] wire_d22_15;
	wire [WIDTH-1:0] wire_d22_16;
	wire [WIDTH-1:0] wire_d22_17;
	wire [WIDTH-1:0] wire_d22_18;
	wire [WIDTH-1:0] wire_d22_19;
	wire [WIDTH-1:0] wire_d22_20;
	wire [WIDTH-1:0] wire_d22_21;
	wire [WIDTH-1:0] wire_d22_22;
	wire [WIDTH-1:0] wire_d22_23;
	wire [WIDTH-1:0] wire_d22_24;
	wire [WIDTH-1:0] wire_d22_25;
	wire [WIDTH-1:0] wire_d22_26;
	wire [WIDTH-1:0] wire_d22_27;
	wire [WIDTH-1:0] wire_d22_28;
	wire [WIDTH-1:0] wire_d22_29;
	wire [WIDTH-1:0] wire_d22_30;
	wire [WIDTH-1:0] wire_d22_31;
	wire [WIDTH-1:0] wire_d22_32;
	wire [WIDTH-1:0] wire_d22_33;
	wire [WIDTH-1:0] wire_d22_34;
	wire [WIDTH-1:0] wire_d22_35;
	wire [WIDTH-1:0] wire_d22_36;
	wire [WIDTH-1:0] wire_d22_37;
	wire [WIDTH-1:0] wire_d22_38;
	wire [WIDTH-1:0] wire_d22_39;
	wire [WIDTH-1:0] wire_d22_40;
	wire [WIDTH-1:0] wire_d22_41;
	wire [WIDTH-1:0] wire_d22_42;
	wire [WIDTH-1:0] wire_d22_43;
	wire [WIDTH-1:0] wire_d22_44;
	wire [WIDTH-1:0] wire_d22_45;
	wire [WIDTH-1:0] wire_d22_46;
	wire [WIDTH-1:0] wire_d22_47;
	wire [WIDTH-1:0] wire_d22_48;
	wire [WIDTH-1:0] wire_d22_49;
	wire [WIDTH-1:0] wire_d22_50;
	wire [WIDTH-1:0] wire_d22_51;
	wire [WIDTH-1:0] wire_d22_52;
	wire [WIDTH-1:0] wire_d22_53;
	wire [WIDTH-1:0] wire_d22_54;
	wire [WIDTH-1:0] wire_d22_55;
	wire [WIDTH-1:0] wire_d22_56;
	wire [WIDTH-1:0] wire_d22_57;
	wire [WIDTH-1:0] wire_d22_58;
	wire [WIDTH-1:0] wire_d22_59;
	wire [WIDTH-1:0] wire_d22_60;
	wire [WIDTH-1:0] wire_d22_61;
	wire [WIDTH-1:0] wire_d22_62;
	wire [WIDTH-1:0] wire_d22_63;
	wire [WIDTH-1:0] wire_d22_64;
	wire [WIDTH-1:0] wire_d22_65;
	wire [WIDTH-1:0] wire_d22_66;
	wire [WIDTH-1:0] wire_d22_67;
	wire [WIDTH-1:0] wire_d22_68;
	wire [WIDTH-1:0] wire_d22_69;
	wire [WIDTH-1:0] wire_d22_70;
	wire [WIDTH-1:0] wire_d22_71;
	wire [WIDTH-1:0] wire_d22_72;
	wire [WIDTH-1:0] wire_d22_73;
	wire [WIDTH-1:0] wire_d22_74;
	wire [WIDTH-1:0] wire_d22_75;
	wire [WIDTH-1:0] wire_d22_76;
	wire [WIDTH-1:0] wire_d22_77;
	wire [WIDTH-1:0] wire_d22_78;
	wire [WIDTH-1:0] wire_d23_0;
	wire [WIDTH-1:0] wire_d23_1;
	wire [WIDTH-1:0] wire_d23_2;
	wire [WIDTH-1:0] wire_d23_3;
	wire [WIDTH-1:0] wire_d23_4;
	wire [WIDTH-1:0] wire_d23_5;
	wire [WIDTH-1:0] wire_d23_6;
	wire [WIDTH-1:0] wire_d23_7;
	wire [WIDTH-1:0] wire_d23_8;
	wire [WIDTH-1:0] wire_d23_9;
	wire [WIDTH-1:0] wire_d23_10;
	wire [WIDTH-1:0] wire_d23_11;
	wire [WIDTH-1:0] wire_d23_12;
	wire [WIDTH-1:0] wire_d23_13;
	wire [WIDTH-1:0] wire_d23_14;
	wire [WIDTH-1:0] wire_d23_15;
	wire [WIDTH-1:0] wire_d23_16;
	wire [WIDTH-1:0] wire_d23_17;
	wire [WIDTH-1:0] wire_d23_18;
	wire [WIDTH-1:0] wire_d23_19;
	wire [WIDTH-1:0] wire_d23_20;
	wire [WIDTH-1:0] wire_d23_21;
	wire [WIDTH-1:0] wire_d23_22;
	wire [WIDTH-1:0] wire_d23_23;
	wire [WIDTH-1:0] wire_d23_24;
	wire [WIDTH-1:0] wire_d23_25;
	wire [WIDTH-1:0] wire_d23_26;
	wire [WIDTH-1:0] wire_d23_27;
	wire [WIDTH-1:0] wire_d23_28;
	wire [WIDTH-1:0] wire_d23_29;
	wire [WIDTH-1:0] wire_d23_30;
	wire [WIDTH-1:0] wire_d23_31;
	wire [WIDTH-1:0] wire_d23_32;
	wire [WIDTH-1:0] wire_d23_33;
	wire [WIDTH-1:0] wire_d23_34;
	wire [WIDTH-1:0] wire_d23_35;
	wire [WIDTH-1:0] wire_d23_36;
	wire [WIDTH-1:0] wire_d23_37;
	wire [WIDTH-1:0] wire_d23_38;
	wire [WIDTH-1:0] wire_d23_39;
	wire [WIDTH-1:0] wire_d23_40;
	wire [WIDTH-1:0] wire_d23_41;
	wire [WIDTH-1:0] wire_d23_42;
	wire [WIDTH-1:0] wire_d23_43;
	wire [WIDTH-1:0] wire_d23_44;
	wire [WIDTH-1:0] wire_d23_45;
	wire [WIDTH-1:0] wire_d23_46;
	wire [WIDTH-1:0] wire_d23_47;
	wire [WIDTH-1:0] wire_d23_48;
	wire [WIDTH-1:0] wire_d23_49;
	wire [WIDTH-1:0] wire_d23_50;
	wire [WIDTH-1:0] wire_d23_51;
	wire [WIDTH-1:0] wire_d23_52;
	wire [WIDTH-1:0] wire_d23_53;
	wire [WIDTH-1:0] wire_d23_54;
	wire [WIDTH-1:0] wire_d23_55;
	wire [WIDTH-1:0] wire_d23_56;
	wire [WIDTH-1:0] wire_d23_57;
	wire [WIDTH-1:0] wire_d23_58;
	wire [WIDTH-1:0] wire_d23_59;
	wire [WIDTH-1:0] wire_d23_60;
	wire [WIDTH-1:0] wire_d23_61;
	wire [WIDTH-1:0] wire_d23_62;
	wire [WIDTH-1:0] wire_d23_63;
	wire [WIDTH-1:0] wire_d23_64;
	wire [WIDTH-1:0] wire_d23_65;
	wire [WIDTH-1:0] wire_d23_66;
	wire [WIDTH-1:0] wire_d23_67;
	wire [WIDTH-1:0] wire_d23_68;
	wire [WIDTH-1:0] wire_d23_69;
	wire [WIDTH-1:0] wire_d23_70;
	wire [WIDTH-1:0] wire_d23_71;
	wire [WIDTH-1:0] wire_d23_72;
	wire [WIDTH-1:0] wire_d23_73;
	wire [WIDTH-1:0] wire_d23_74;
	wire [WIDTH-1:0] wire_d23_75;
	wire [WIDTH-1:0] wire_d23_76;
	wire [WIDTH-1:0] wire_d23_77;
	wire [WIDTH-1:0] wire_d23_78;
	wire [WIDTH-1:0] wire_d24_0;
	wire [WIDTH-1:0] wire_d24_1;
	wire [WIDTH-1:0] wire_d24_2;
	wire [WIDTH-1:0] wire_d24_3;
	wire [WIDTH-1:0] wire_d24_4;
	wire [WIDTH-1:0] wire_d24_5;
	wire [WIDTH-1:0] wire_d24_6;
	wire [WIDTH-1:0] wire_d24_7;
	wire [WIDTH-1:0] wire_d24_8;
	wire [WIDTH-1:0] wire_d24_9;
	wire [WIDTH-1:0] wire_d24_10;
	wire [WIDTH-1:0] wire_d24_11;
	wire [WIDTH-1:0] wire_d24_12;
	wire [WIDTH-1:0] wire_d24_13;
	wire [WIDTH-1:0] wire_d24_14;
	wire [WIDTH-1:0] wire_d24_15;
	wire [WIDTH-1:0] wire_d24_16;
	wire [WIDTH-1:0] wire_d24_17;
	wire [WIDTH-1:0] wire_d24_18;
	wire [WIDTH-1:0] wire_d24_19;
	wire [WIDTH-1:0] wire_d24_20;
	wire [WIDTH-1:0] wire_d24_21;
	wire [WIDTH-1:0] wire_d24_22;
	wire [WIDTH-1:0] wire_d24_23;
	wire [WIDTH-1:0] wire_d24_24;
	wire [WIDTH-1:0] wire_d24_25;
	wire [WIDTH-1:0] wire_d24_26;
	wire [WIDTH-1:0] wire_d24_27;
	wire [WIDTH-1:0] wire_d24_28;
	wire [WIDTH-1:0] wire_d24_29;
	wire [WIDTH-1:0] wire_d24_30;
	wire [WIDTH-1:0] wire_d24_31;
	wire [WIDTH-1:0] wire_d24_32;
	wire [WIDTH-1:0] wire_d24_33;
	wire [WIDTH-1:0] wire_d24_34;
	wire [WIDTH-1:0] wire_d24_35;
	wire [WIDTH-1:0] wire_d24_36;
	wire [WIDTH-1:0] wire_d24_37;
	wire [WIDTH-1:0] wire_d24_38;
	wire [WIDTH-1:0] wire_d24_39;
	wire [WIDTH-1:0] wire_d24_40;
	wire [WIDTH-1:0] wire_d24_41;
	wire [WIDTH-1:0] wire_d24_42;
	wire [WIDTH-1:0] wire_d24_43;
	wire [WIDTH-1:0] wire_d24_44;
	wire [WIDTH-1:0] wire_d24_45;
	wire [WIDTH-1:0] wire_d24_46;
	wire [WIDTH-1:0] wire_d24_47;
	wire [WIDTH-1:0] wire_d24_48;
	wire [WIDTH-1:0] wire_d24_49;
	wire [WIDTH-1:0] wire_d24_50;
	wire [WIDTH-1:0] wire_d24_51;
	wire [WIDTH-1:0] wire_d24_52;
	wire [WIDTH-1:0] wire_d24_53;
	wire [WIDTH-1:0] wire_d24_54;
	wire [WIDTH-1:0] wire_d24_55;
	wire [WIDTH-1:0] wire_d24_56;
	wire [WIDTH-1:0] wire_d24_57;
	wire [WIDTH-1:0] wire_d24_58;
	wire [WIDTH-1:0] wire_d24_59;
	wire [WIDTH-1:0] wire_d24_60;
	wire [WIDTH-1:0] wire_d24_61;
	wire [WIDTH-1:0] wire_d24_62;
	wire [WIDTH-1:0] wire_d24_63;
	wire [WIDTH-1:0] wire_d24_64;
	wire [WIDTH-1:0] wire_d24_65;
	wire [WIDTH-1:0] wire_d24_66;
	wire [WIDTH-1:0] wire_d24_67;
	wire [WIDTH-1:0] wire_d24_68;
	wire [WIDTH-1:0] wire_d24_69;
	wire [WIDTH-1:0] wire_d24_70;
	wire [WIDTH-1:0] wire_d24_71;
	wire [WIDTH-1:0] wire_d24_72;
	wire [WIDTH-1:0] wire_d24_73;
	wire [WIDTH-1:0] wire_d24_74;
	wire [WIDTH-1:0] wire_d24_75;
	wire [WIDTH-1:0] wire_d24_76;
	wire [WIDTH-1:0] wire_d24_77;
	wire [WIDTH-1:0] wire_d24_78;
	wire [WIDTH-1:0] wire_d25_0;
	wire [WIDTH-1:0] wire_d25_1;
	wire [WIDTH-1:0] wire_d25_2;
	wire [WIDTH-1:0] wire_d25_3;
	wire [WIDTH-1:0] wire_d25_4;
	wire [WIDTH-1:0] wire_d25_5;
	wire [WIDTH-1:0] wire_d25_6;
	wire [WIDTH-1:0] wire_d25_7;
	wire [WIDTH-1:0] wire_d25_8;
	wire [WIDTH-1:0] wire_d25_9;
	wire [WIDTH-1:0] wire_d25_10;
	wire [WIDTH-1:0] wire_d25_11;
	wire [WIDTH-1:0] wire_d25_12;
	wire [WIDTH-1:0] wire_d25_13;
	wire [WIDTH-1:0] wire_d25_14;
	wire [WIDTH-1:0] wire_d25_15;
	wire [WIDTH-1:0] wire_d25_16;
	wire [WIDTH-1:0] wire_d25_17;
	wire [WIDTH-1:0] wire_d25_18;
	wire [WIDTH-1:0] wire_d25_19;
	wire [WIDTH-1:0] wire_d25_20;
	wire [WIDTH-1:0] wire_d25_21;
	wire [WIDTH-1:0] wire_d25_22;
	wire [WIDTH-1:0] wire_d25_23;
	wire [WIDTH-1:0] wire_d25_24;
	wire [WIDTH-1:0] wire_d25_25;
	wire [WIDTH-1:0] wire_d25_26;
	wire [WIDTH-1:0] wire_d25_27;
	wire [WIDTH-1:0] wire_d25_28;
	wire [WIDTH-1:0] wire_d25_29;
	wire [WIDTH-1:0] wire_d25_30;
	wire [WIDTH-1:0] wire_d25_31;
	wire [WIDTH-1:0] wire_d25_32;
	wire [WIDTH-1:0] wire_d25_33;
	wire [WIDTH-1:0] wire_d25_34;
	wire [WIDTH-1:0] wire_d25_35;
	wire [WIDTH-1:0] wire_d25_36;
	wire [WIDTH-1:0] wire_d25_37;
	wire [WIDTH-1:0] wire_d25_38;
	wire [WIDTH-1:0] wire_d25_39;
	wire [WIDTH-1:0] wire_d25_40;
	wire [WIDTH-1:0] wire_d25_41;
	wire [WIDTH-1:0] wire_d25_42;
	wire [WIDTH-1:0] wire_d25_43;
	wire [WIDTH-1:0] wire_d25_44;
	wire [WIDTH-1:0] wire_d25_45;
	wire [WIDTH-1:0] wire_d25_46;
	wire [WIDTH-1:0] wire_d25_47;
	wire [WIDTH-1:0] wire_d25_48;
	wire [WIDTH-1:0] wire_d25_49;
	wire [WIDTH-1:0] wire_d25_50;
	wire [WIDTH-1:0] wire_d25_51;
	wire [WIDTH-1:0] wire_d25_52;
	wire [WIDTH-1:0] wire_d25_53;
	wire [WIDTH-1:0] wire_d25_54;
	wire [WIDTH-1:0] wire_d25_55;
	wire [WIDTH-1:0] wire_d25_56;
	wire [WIDTH-1:0] wire_d25_57;
	wire [WIDTH-1:0] wire_d25_58;
	wire [WIDTH-1:0] wire_d25_59;
	wire [WIDTH-1:0] wire_d25_60;
	wire [WIDTH-1:0] wire_d25_61;
	wire [WIDTH-1:0] wire_d25_62;
	wire [WIDTH-1:0] wire_d25_63;
	wire [WIDTH-1:0] wire_d25_64;
	wire [WIDTH-1:0] wire_d25_65;
	wire [WIDTH-1:0] wire_d25_66;
	wire [WIDTH-1:0] wire_d25_67;
	wire [WIDTH-1:0] wire_d25_68;
	wire [WIDTH-1:0] wire_d25_69;
	wire [WIDTH-1:0] wire_d25_70;
	wire [WIDTH-1:0] wire_d25_71;
	wire [WIDTH-1:0] wire_d25_72;
	wire [WIDTH-1:0] wire_d25_73;
	wire [WIDTH-1:0] wire_d25_74;
	wire [WIDTH-1:0] wire_d25_75;
	wire [WIDTH-1:0] wire_d25_76;
	wire [WIDTH-1:0] wire_d25_77;
	wire [WIDTH-1:0] wire_d25_78;
	wire [WIDTH-1:0] wire_d26_0;
	wire [WIDTH-1:0] wire_d26_1;
	wire [WIDTH-1:0] wire_d26_2;
	wire [WIDTH-1:0] wire_d26_3;
	wire [WIDTH-1:0] wire_d26_4;
	wire [WIDTH-1:0] wire_d26_5;
	wire [WIDTH-1:0] wire_d26_6;
	wire [WIDTH-1:0] wire_d26_7;
	wire [WIDTH-1:0] wire_d26_8;
	wire [WIDTH-1:0] wire_d26_9;
	wire [WIDTH-1:0] wire_d26_10;
	wire [WIDTH-1:0] wire_d26_11;
	wire [WIDTH-1:0] wire_d26_12;
	wire [WIDTH-1:0] wire_d26_13;
	wire [WIDTH-1:0] wire_d26_14;
	wire [WIDTH-1:0] wire_d26_15;
	wire [WIDTH-1:0] wire_d26_16;
	wire [WIDTH-1:0] wire_d26_17;
	wire [WIDTH-1:0] wire_d26_18;
	wire [WIDTH-1:0] wire_d26_19;
	wire [WIDTH-1:0] wire_d26_20;
	wire [WIDTH-1:0] wire_d26_21;
	wire [WIDTH-1:0] wire_d26_22;
	wire [WIDTH-1:0] wire_d26_23;
	wire [WIDTH-1:0] wire_d26_24;
	wire [WIDTH-1:0] wire_d26_25;
	wire [WIDTH-1:0] wire_d26_26;
	wire [WIDTH-1:0] wire_d26_27;
	wire [WIDTH-1:0] wire_d26_28;
	wire [WIDTH-1:0] wire_d26_29;
	wire [WIDTH-1:0] wire_d26_30;
	wire [WIDTH-1:0] wire_d26_31;
	wire [WIDTH-1:0] wire_d26_32;
	wire [WIDTH-1:0] wire_d26_33;
	wire [WIDTH-1:0] wire_d26_34;
	wire [WIDTH-1:0] wire_d26_35;
	wire [WIDTH-1:0] wire_d26_36;
	wire [WIDTH-1:0] wire_d26_37;
	wire [WIDTH-1:0] wire_d26_38;
	wire [WIDTH-1:0] wire_d26_39;
	wire [WIDTH-1:0] wire_d26_40;
	wire [WIDTH-1:0] wire_d26_41;
	wire [WIDTH-1:0] wire_d26_42;
	wire [WIDTH-1:0] wire_d26_43;
	wire [WIDTH-1:0] wire_d26_44;
	wire [WIDTH-1:0] wire_d26_45;
	wire [WIDTH-1:0] wire_d26_46;
	wire [WIDTH-1:0] wire_d26_47;
	wire [WIDTH-1:0] wire_d26_48;
	wire [WIDTH-1:0] wire_d26_49;
	wire [WIDTH-1:0] wire_d26_50;
	wire [WIDTH-1:0] wire_d26_51;
	wire [WIDTH-1:0] wire_d26_52;
	wire [WIDTH-1:0] wire_d26_53;
	wire [WIDTH-1:0] wire_d26_54;
	wire [WIDTH-1:0] wire_d26_55;
	wire [WIDTH-1:0] wire_d26_56;
	wire [WIDTH-1:0] wire_d26_57;
	wire [WIDTH-1:0] wire_d26_58;
	wire [WIDTH-1:0] wire_d26_59;
	wire [WIDTH-1:0] wire_d26_60;
	wire [WIDTH-1:0] wire_d26_61;
	wire [WIDTH-1:0] wire_d26_62;
	wire [WIDTH-1:0] wire_d26_63;
	wire [WIDTH-1:0] wire_d26_64;
	wire [WIDTH-1:0] wire_d26_65;
	wire [WIDTH-1:0] wire_d26_66;
	wire [WIDTH-1:0] wire_d26_67;
	wire [WIDTH-1:0] wire_d26_68;
	wire [WIDTH-1:0] wire_d26_69;
	wire [WIDTH-1:0] wire_d26_70;
	wire [WIDTH-1:0] wire_d26_71;
	wire [WIDTH-1:0] wire_d26_72;
	wire [WIDTH-1:0] wire_d26_73;
	wire [WIDTH-1:0] wire_d26_74;
	wire [WIDTH-1:0] wire_d26_75;
	wire [WIDTH-1:0] wire_d26_76;
	wire [WIDTH-1:0] wire_d26_77;
	wire [WIDTH-1:0] wire_d26_78;
	wire [WIDTH-1:0] wire_d27_0;
	wire [WIDTH-1:0] wire_d27_1;
	wire [WIDTH-1:0] wire_d27_2;
	wire [WIDTH-1:0] wire_d27_3;
	wire [WIDTH-1:0] wire_d27_4;
	wire [WIDTH-1:0] wire_d27_5;
	wire [WIDTH-1:0] wire_d27_6;
	wire [WIDTH-1:0] wire_d27_7;
	wire [WIDTH-1:0] wire_d27_8;
	wire [WIDTH-1:0] wire_d27_9;
	wire [WIDTH-1:0] wire_d27_10;
	wire [WIDTH-1:0] wire_d27_11;
	wire [WIDTH-1:0] wire_d27_12;
	wire [WIDTH-1:0] wire_d27_13;
	wire [WIDTH-1:0] wire_d27_14;
	wire [WIDTH-1:0] wire_d27_15;
	wire [WIDTH-1:0] wire_d27_16;
	wire [WIDTH-1:0] wire_d27_17;
	wire [WIDTH-1:0] wire_d27_18;
	wire [WIDTH-1:0] wire_d27_19;
	wire [WIDTH-1:0] wire_d27_20;
	wire [WIDTH-1:0] wire_d27_21;
	wire [WIDTH-1:0] wire_d27_22;
	wire [WIDTH-1:0] wire_d27_23;
	wire [WIDTH-1:0] wire_d27_24;
	wire [WIDTH-1:0] wire_d27_25;
	wire [WIDTH-1:0] wire_d27_26;
	wire [WIDTH-1:0] wire_d27_27;
	wire [WIDTH-1:0] wire_d27_28;
	wire [WIDTH-1:0] wire_d27_29;
	wire [WIDTH-1:0] wire_d27_30;
	wire [WIDTH-1:0] wire_d27_31;
	wire [WIDTH-1:0] wire_d27_32;
	wire [WIDTH-1:0] wire_d27_33;
	wire [WIDTH-1:0] wire_d27_34;
	wire [WIDTH-1:0] wire_d27_35;
	wire [WIDTH-1:0] wire_d27_36;
	wire [WIDTH-1:0] wire_d27_37;
	wire [WIDTH-1:0] wire_d27_38;
	wire [WIDTH-1:0] wire_d27_39;
	wire [WIDTH-1:0] wire_d27_40;
	wire [WIDTH-1:0] wire_d27_41;
	wire [WIDTH-1:0] wire_d27_42;
	wire [WIDTH-1:0] wire_d27_43;
	wire [WIDTH-1:0] wire_d27_44;
	wire [WIDTH-1:0] wire_d27_45;
	wire [WIDTH-1:0] wire_d27_46;
	wire [WIDTH-1:0] wire_d27_47;
	wire [WIDTH-1:0] wire_d27_48;
	wire [WIDTH-1:0] wire_d27_49;
	wire [WIDTH-1:0] wire_d27_50;
	wire [WIDTH-1:0] wire_d27_51;
	wire [WIDTH-1:0] wire_d27_52;
	wire [WIDTH-1:0] wire_d27_53;
	wire [WIDTH-1:0] wire_d27_54;
	wire [WIDTH-1:0] wire_d27_55;
	wire [WIDTH-1:0] wire_d27_56;
	wire [WIDTH-1:0] wire_d27_57;
	wire [WIDTH-1:0] wire_d27_58;
	wire [WIDTH-1:0] wire_d27_59;
	wire [WIDTH-1:0] wire_d27_60;
	wire [WIDTH-1:0] wire_d27_61;
	wire [WIDTH-1:0] wire_d27_62;
	wire [WIDTH-1:0] wire_d27_63;
	wire [WIDTH-1:0] wire_d27_64;
	wire [WIDTH-1:0] wire_d27_65;
	wire [WIDTH-1:0] wire_d27_66;
	wire [WIDTH-1:0] wire_d27_67;
	wire [WIDTH-1:0] wire_d27_68;
	wire [WIDTH-1:0] wire_d27_69;
	wire [WIDTH-1:0] wire_d27_70;
	wire [WIDTH-1:0] wire_d27_71;
	wire [WIDTH-1:0] wire_d27_72;
	wire [WIDTH-1:0] wire_d27_73;
	wire [WIDTH-1:0] wire_d27_74;
	wire [WIDTH-1:0] wire_d27_75;
	wire [WIDTH-1:0] wire_d27_76;
	wire [WIDTH-1:0] wire_d27_77;
	wire [WIDTH-1:0] wire_d27_78;
	wire [WIDTH-1:0] wire_d28_0;
	wire [WIDTH-1:0] wire_d28_1;
	wire [WIDTH-1:0] wire_d28_2;
	wire [WIDTH-1:0] wire_d28_3;
	wire [WIDTH-1:0] wire_d28_4;
	wire [WIDTH-1:0] wire_d28_5;
	wire [WIDTH-1:0] wire_d28_6;
	wire [WIDTH-1:0] wire_d28_7;
	wire [WIDTH-1:0] wire_d28_8;
	wire [WIDTH-1:0] wire_d28_9;
	wire [WIDTH-1:0] wire_d28_10;
	wire [WIDTH-1:0] wire_d28_11;
	wire [WIDTH-1:0] wire_d28_12;
	wire [WIDTH-1:0] wire_d28_13;
	wire [WIDTH-1:0] wire_d28_14;
	wire [WIDTH-1:0] wire_d28_15;
	wire [WIDTH-1:0] wire_d28_16;
	wire [WIDTH-1:0] wire_d28_17;
	wire [WIDTH-1:0] wire_d28_18;
	wire [WIDTH-1:0] wire_d28_19;
	wire [WIDTH-1:0] wire_d28_20;
	wire [WIDTH-1:0] wire_d28_21;
	wire [WIDTH-1:0] wire_d28_22;
	wire [WIDTH-1:0] wire_d28_23;
	wire [WIDTH-1:0] wire_d28_24;
	wire [WIDTH-1:0] wire_d28_25;
	wire [WIDTH-1:0] wire_d28_26;
	wire [WIDTH-1:0] wire_d28_27;
	wire [WIDTH-1:0] wire_d28_28;
	wire [WIDTH-1:0] wire_d28_29;
	wire [WIDTH-1:0] wire_d28_30;
	wire [WIDTH-1:0] wire_d28_31;
	wire [WIDTH-1:0] wire_d28_32;
	wire [WIDTH-1:0] wire_d28_33;
	wire [WIDTH-1:0] wire_d28_34;
	wire [WIDTH-1:0] wire_d28_35;
	wire [WIDTH-1:0] wire_d28_36;
	wire [WIDTH-1:0] wire_d28_37;
	wire [WIDTH-1:0] wire_d28_38;
	wire [WIDTH-1:0] wire_d28_39;
	wire [WIDTH-1:0] wire_d28_40;
	wire [WIDTH-1:0] wire_d28_41;
	wire [WIDTH-1:0] wire_d28_42;
	wire [WIDTH-1:0] wire_d28_43;
	wire [WIDTH-1:0] wire_d28_44;
	wire [WIDTH-1:0] wire_d28_45;
	wire [WIDTH-1:0] wire_d28_46;
	wire [WIDTH-1:0] wire_d28_47;
	wire [WIDTH-1:0] wire_d28_48;
	wire [WIDTH-1:0] wire_d28_49;
	wire [WIDTH-1:0] wire_d28_50;
	wire [WIDTH-1:0] wire_d28_51;
	wire [WIDTH-1:0] wire_d28_52;
	wire [WIDTH-1:0] wire_d28_53;
	wire [WIDTH-1:0] wire_d28_54;
	wire [WIDTH-1:0] wire_d28_55;
	wire [WIDTH-1:0] wire_d28_56;
	wire [WIDTH-1:0] wire_d28_57;
	wire [WIDTH-1:0] wire_d28_58;
	wire [WIDTH-1:0] wire_d28_59;
	wire [WIDTH-1:0] wire_d28_60;
	wire [WIDTH-1:0] wire_d28_61;
	wire [WIDTH-1:0] wire_d28_62;
	wire [WIDTH-1:0] wire_d28_63;
	wire [WIDTH-1:0] wire_d28_64;
	wire [WIDTH-1:0] wire_d28_65;
	wire [WIDTH-1:0] wire_d28_66;
	wire [WIDTH-1:0] wire_d28_67;
	wire [WIDTH-1:0] wire_d28_68;
	wire [WIDTH-1:0] wire_d28_69;
	wire [WIDTH-1:0] wire_d28_70;
	wire [WIDTH-1:0] wire_d28_71;
	wire [WIDTH-1:0] wire_d28_72;
	wire [WIDTH-1:0] wire_d28_73;
	wire [WIDTH-1:0] wire_d28_74;
	wire [WIDTH-1:0] wire_d28_75;
	wire [WIDTH-1:0] wire_d28_76;
	wire [WIDTH-1:0] wire_d28_77;
	wire [WIDTH-1:0] wire_d28_78;
	wire [WIDTH-1:0] wire_d29_0;
	wire [WIDTH-1:0] wire_d29_1;
	wire [WIDTH-1:0] wire_d29_2;
	wire [WIDTH-1:0] wire_d29_3;
	wire [WIDTH-1:0] wire_d29_4;
	wire [WIDTH-1:0] wire_d29_5;
	wire [WIDTH-1:0] wire_d29_6;
	wire [WIDTH-1:0] wire_d29_7;
	wire [WIDTH-1:0] wire_d29_8;
	wire [WIDTH-1:0] wire_d29_9;
	wire [WIDTH-1:0] wire_d29_10;
	wire [WIDTH-1:0] wire_d29_11;
	wire [WIDTH-1:0] wire_d29_12;
	wire [WIDTH-1:0] wire_d29_13;
	wire [WIDTH-1:0] wire_d29_14;
	wire [WIDTH-1:0] wire_d29_15;
	wire [WIDTH-1:0] wire_d29_16;
	wire [WIDTH-1:0] wire_d29_17;
	wire [WIDTH-1:0] wire_d29_18;
	wire [WIDTH-1:0] wire_d29_19;
	wire [WIDTH-1:0] wire_d29_20;
	wire [WIDTH-1:0] wire_d29_21;
	wire [WIDTH-1:0] wire_d29_22;
	wire [WIDTH-1:0] wire_d29_23;
	wire [WIDTH-1:0] wire_d29_24;
	wire [WIDTH-1:0] wire_d29_25;
	wire [WIDTH-1:0] wire_d29_26;
	wire [WIDTH-1:0] wire_d29_27;
	wire [WIDTH-1:0] wire_d29_28;
	wire [WIDTH-1:0] wire_d29_29;
	wire [WIDTH-1:0] wire_d29_30;
	wire [WIDTH-1:0] wire_d29_31;
	wire [WIDTH-1:0] wire_d29_32;
	wire [WIDTH-1:0] wire_d29_33;
	wire [WIDTH-1:0] wire_d29_34;
	wire [WIDTH-1:0] wire_d29_35;
	wire [WIDTH-1:0] wire_d29_36;
	wire [WIDTH-1:0] wire_d29_37;
	wire [WIDTH-1:0] wire_d29_38;
	wire [WIDTH-1:0] wire_d29_39;
	wire [WIDTH-1:0] wire_d29_40;
	wire [WIDTH-1:0] wire_d29_41;
	wire [WIDTH-1:0] wire_d29_42;
	wire [WIDTH-1:0] wire_d29_43;
	wire [WIDTH-1:0] wire_d29_44;
	wire [WIDTH-1:0] wire_d29_45;
	wire [WIDTH-1:0] wire_d29_46;
	wire [WIDTH-1:0] wire_d29_47;
	wire [WIDTH-1:0] wire_d29_48;
	wire [WIDTH-1:0] wire_d29_49;
	wire [WIDTH-1:0] wire_d29_50;
	wire [WIDTH-1:0] wire_d29_51;
	wire [WIDTH-1:0] wire_d29_52;
	wire [WIDTH-1:0] wire_d29_53;
	wire [WIDTH-1:0] wire_d29_54;
	wire [WIDTH-1:0] wire_d29_55;
	wire [WIDTH-1:0] wire_d29_56;
	wire [WIDTH-1:0] wire_d29_57;
	wire [WIDTH-1:0] wire_d29_58;
	wire [WIDTH-1:0] wire_d29_59;
	wire [WIDTH-1:0] wire_d29_60;
	wire [WIDTH-1:0] wire_d29_61;
	wire [WIDTH-1:0] wire_d29_62;
	wire [WIDTH-1:0] wire_d29_63;
	wire [WIDTH-1:0] wire_d29_64;
	wire [WIDTH-1:0] wire_d29_65;
	wire [WIDTH-1:0] wire_d29_66;
	wire [WIDTH-1:0] wire_d29_67;
	wire [WIDTH-1:0] wire_d29_68;
	wire [WIDTH-1:0] wire_d29_69;
	wire [WIDTH-1:0] wire_d29_70;
	wire [WIDTH-1:0] wire_d29_71;
	wire [WIDTH-1:0] wire_d29_72;
	wire [WIDTH-1:0] wire_d29_73;
	wire [WIDTH-1:0] wire_d29_74;
	wire [WIDTH-1:0] wire_d29_75;
	wire [WIDTH-1:0] wire_d29_76;
	wire [WIDTH-1:0] wire_d29_77;
	wire [WIDTH-1:0] wire_d29_78;
	wire [WIDTH-1:0] wire_d30_0;
	wire [WIDTH-1:0] wire_d30_1;
	wire [WIDTH-1:0] wire_d30_2;
	wire [WIDTH-1:0] wire_d30_3;
	wire [WIDTH-1:0] wire_d30_4;
	wire [WIDTH-1:0] wire_d30_5;
	wire [WIDTH-1:0] wire_d30_6;
	wire [WIDTH-1:0] wire_d30_7;
	wire [WIDTH-1:0] wire_d30_8;
	wire [WIDTH-1:0] wire_d30_9;
	wire [WIDTH-1:0] wire_d30_10;
	wire [WIDTH-1:0] wire_d30_11;
	wire [WIDTH-1:0] wire_d30_12;
	wire [WIDTH-1:0] wire_d30_13;
	wire [WIDTH-1:0] wire_d30_14;
	wire [WIDTH-1:0] wire_d30_15;
	wire [WIDTH-1:0] wire_d30_16;
	wire [WIDTH-1:0] wire_d30_17;
	wire [WIDTH-1:0] wire_d30_18;
	wire [WIDTH-1:0] wire_d30_19;
	wire [WIDTH-1:0] wire_d30_20;
	wire [WIDTH-1:0] wire_d30_21;
	wire [WIDTH-1:0] wire_d30_22;
	wire [WIDTH-1:0] wire_d30_23;
	wire [WIDTH-1:0] wire_d30_24;
	wire [WIDTH-1:0] wire_d30_25;
	wire [WIDTH-1:0] wire_d30_26;
	wire [WIDTH-1:0] wire_d30_27;
	wire [WIDTH-1:0] wire_d30_28;
	wire [WIDTH-1:0] wire_d30_29;
	wire [WIDTH-1:0] wire_d30_30;
	wire [WIDTH-1:0] wire_d30_31;
	wire [WIDTH-1:0] wire_d30_32;
	wire [WIDTH-1:0] wire_d30_33;
	wire [WIDTH-1:0] wire_d30_34;
	wire [WIDTH-1:0] wire_d30_35;
	wire [WIDTH-1:0] wire_d30_36;
	wire [WIDTH-1:0] wire_d30_37;
	wire [WIDTH-1:0] wire_d30_38;
	wire [WIDTH-1:0] wire_d30_39;
	wire [WIDTH-1:0] wire_d30_40;
	wire [WIDTH-1:0] wire_d30_41;
	wire [WIDTH-1:0] wire_d30_42;
	wire [WIDTH-1:0] wire_d30_43;
	wire [WIDTH-1:0] wire_d30_44;
	wire [WIDTH-1:0] wire_d30_45;
	wire [WIDTH-1:0] wire_d30_46;
	wire [WIDTH-1:0] wire_d30_47;
	wire [WIDTH-1:0] wire_d30_48;
	wire [WIDTH-1:0] wire_d30_49;
	wire [WIDTH-1:0] wire_d30_50;
	wire [WIDTH-1:0] wire_d30_51;
	wire [WIDTH-1:0] wire_d30_52;
	wire [WIDTH-1:0] wire_d30_53;
	wire [WIDTH-1:0] wire_d30_54;
	wire [WIDTH-1:0] wire_d30_55;
	wire [WIDTH-1:0] wire_d30_56;
	wire [WIDTH-1:0] wire_d30_57;
	wire [WIDTH-1:0] wire_d30_58;
	wire [WIDTH-1:0] wire_d30_59;
	wire [WIDTH-1:0] wire_d30_60;
	wire [WIDTH-1:0] wire_d30_61;
	wire [WIDTH-1:0] wire_d30_62;
	wire [WIDTH-1:0] wire_d30_63;
	wire [WIDTH-1:0] wire_d30_64;
	wire [WIDTH-1:0] wire_d30_65;
	wire [WIDTH-1:0] wire_d30_66;
	wire [WIDTH-1:0] wire_d30_67;
	wire [WIDTH-1:0] wire_d30_68;
	wire [WIDTH-1:0] wire_d30_69;
	wire [WIDTH-1:0] wire_d30_70;
	wire [WIDTH-1:0] wire_d30_71;
	wire [WIDTH-1:0] wire_d30_72;
	wire [WIDTH-1:0] wire_d30_73;
	wire [WIDTH-1:0] wire_d30_74;
	wire [WIDTH-1:0] wire_d30_75;
	wire [WIDTH-1:0] wire_d30_76;
	wire [WIDTH-1:0] wire_d30_77;
	wire [WIDTH-1:0] wire_d30_78;
	wire [WIDTH-1:0] wire_d31_0;
	wire [WIDTH-1:0] wire_d31_1;
	wire [WIDTH-1:0] wire_d31_2;
	wire [WIDTH-1:0] wire_d31_3;
	wire [WIDTH-1:0] wire_d31_4;
	wire [WIDTH-1:0] wire_d31_5;
	wire [WIDTH-1:0] wire_d31_6;
	wire [WIDTH-1:0] wire_d31_7;
	wire [WIDTH-1:0] wire_d31_8;
	wire [WIDTH-1:0] wire_d31_9;
	wire [WIDTH-1:0] wire_d31_10;
	wire [WIDTH-1:0] wire_d31_11;
	wire [WIDTH-1:0] wire_d31_12;
	wire [WIDTH-1:0] wire_d31_13;
	wire [WIDTH-1:0] wire_d31_14;
	wire [WIDTH-1:0] wire_d31_15;
	wire [WIDTH-1:0] wire_d31_16;
	wire [WIDTH-1:0] wire_d31_17;
	wire [WIDTH-1:0] wire_d31_18;
	wire [WIDTH-1:0] wire_d31_19;
	wire [WIDTH-1:0] wire_d31_20;
	wire [WIDTH-1:0] wire_d31_21;
	wire [WIDTH-1:0] wire_d31_22;
	wire [WIDTH-1:0] wire_d31_23;
	wire [WIDTH-1:0] wire_d31_24;
	wire [WIDTH-1:0] wire_d31_25;
	wire [WIDTH-1:0] wire_d31_26;
	wire [WIDTH-1:0] wire_d31_27;
	wire [WIDTH-1:0] wire_d31_28;
	wire [WIDTH-1:0] wire_d31_29;
	wire [WIDTH-1:0] wire_d31_30;
	wire [WIDTH-1:0] wire_d31_31;
	wire [WIDTH-1:0] wire_d31_32;
	wire [WIDTH-1:0] wire_d31_33;
	wire [WIDTH-1:0] wire_d31_34;
	wire [WIDTH-1:0] wire_d31_35;
	wire [WIDTH-1:0] wire_d31_36;
	wire [WIDTH-1:0] wire_d31_37;
	wire [WIDTH-1:0] wire_d31_38;
	wire [WIDTH-1:0] wire_d31_39;
	wire [WIDTH-1:0] wire_d31_40;
	wire [WIDTH-1:0] wire_d31_41;
	wire [WIDTH-1:0] wire_d31_42;
	wire [WIDTH-1:0] wire_d31_43;
	wire [WIDTH-1:0] wire_d31_44;
	wire [WIDTH-1:0] wire_d31_45;
	wire [WIDTH-1:0] wire_d31_46;
	wire [WIDTH-1:0] wire_d31_47;
	wire [WIDTH-1:0] wire_d31_48;
	wire [WIDTH-1:0] wire_d31_49;
	wire [WIDTH-1:0] wire_d31_50;
	wire [WIDTH-1:0] wire_d31_51;
	wire [WIDTH-1:0] wire_d31_52;
	wire [WIDTH-1:0] wire_d31_53;
	wire [WIDTH-1:0] wire_d31_54;
	wire [WIDTH-1:0] wire_d31_55;
	wire [WIDTH-1:0] wire_d31_56;
	wire [WIDTH-1:0] wire_d31_57;
	wire [WIDTH-1:0] wire_d31_58;
	wire [WIDTH-1:0] wire_d31_59;
	wire [WIDTH-1:0] wire_d31_60;
	wire [WIDTH-1:0] wire_d31_61;
	wire [WIDTH-1:0] wire_d31_62;
	wire [WIDTH-1:0] wire_d31_63;
	wire [WIDTH-1:0] wire_d31_64;
	wire [WIDTH-1:0] wire_d31_65;
	wire [WIDTH-1:0] wire_d31_66;
	wire [WIDTH-1:0] wire_d31_67;
	wire [WIDTH-1:0] wire_d31_68;
	wire [WIDTH-1:0] wire_d31_69;
	wire [WIDTH-1:0] wire_d31_70;
	wire [WIDTH-1:0] wire_d31_71;
	wire [WIDTH-1:0] wire_d31_72;
	wire [WIDTH-1:0] wire_d31_73;
	wire [WIDTH-1:0] wire_d31_74;
	wire [WIDTH-1:0] wire_d31_75;
	wire [WIDTH-1:0] wire_d31_76;
	wire [WIDTH-1:0] wire_d31_77;
	wire [WIDTH-1:0] wire_d31_78;
	wire [WIDTH-1:0] wire_d32_0;
	wire [WIDTH-1:0] wire_d32_1;
	wire [WIDTH-1:0] wire_d32_2;
	wire [WIDTH-1:0] wire_d32_3;
	wire [WIDTH-1:0] wire_d32_4;
	wire [WIDTH-1:0] wire_d32_5;
	wire [WIDTH-1:0] wire_d32_6;
	wire [WIDTH-1:0] wire_d32_7;
	wire [WIDTH-1:0] wire_d32_8;
	wire [WIDTH-1:0] wire_d32_9;
	wire [WIDTH-1:0] wire_d32_10;
	wire [WIDTH-1:0] wire_d32_11;
	wire [WIDTH-1:0] wire_d32_12;
	wire [WIDTH-1:0] wire_d32_13;
	wire [WIDTH-1:0] wire_d32_14;
	wire [WIDTH-1:0] wire_d32_15;
	wire [WIDTH-1:0] wire_d32_16;
	wire [WIDTH-1:0] wire_d32_17;
	wire [WIDTH-1:0] wire_d32_18;
	wire [WIDTH-1:0] wire_d32_19;
	wire [WIDTH-1:0] wire_d32_20;
	wire [WIDTH-1:0] wire_d32_21;
	wire [WIDTH-1:0] wire_d32_22;
	wire [WIDTH-1:0] wire_d32_23;
	wire [WIDTH-1:0] wire_d32_24;
	wire [WIDTH-1:0] wire_d32_25;
	wire [WIDTH-1:0] wire_d32_26;
	wire [WIDTH-1:0] wire_d32_27;
	wire [WIDTH-1:0] wire_d32_28;
	wire [WIDTH-1:0] wire_d32_29;
	wire [WIDTH-1:0] wire_d32_30;
	wire [WIDTH-1:0] wire_d32_31;
	wire [WIDTH-1:0] wire_d32_32;
	wire [WIDTH-1:0] wire_d32_33;
	wire [WIDTH-1:0] wire_d32_34;
	wire [WIDTH-1:0] wire_d32_35;
	wire [WIDTH-1:0] wire_d32_36;
	wire [WIDTH-1:0] wire_d32_37;
	wire [WIDTH-1:0] wire_d32_38;
	wire [WIDTH-1:0] wire_d32_39;
	wire [WIDTH-1:0] wire_d32_40;
	wire [WIDTH-1:0] wire_d32_41;
	wire [WIDTH-1:0] wire_d32_42;
	wire [WIDTH-1:0] wire_d32_43;
	wire [WIDTH-1:0] wire_d32_44;
	wire [WIDTH-1:0] wire_d32_45;
	wire [WIDTH-1:0] wire_d32_46;
	wire [WIDTH-1:0] wire_d32_47;
	wire [WIDTH-1:0] wire_d32_48;
	wire [WIDTH-1:0] wire_d32_49;
	wire [WIDTH-1:0] wire_d32_50;
	wire [WIDTH-1:0] wire_d32_51;
	wire [WIDTH-1:0] wire_d32_52;
	wire [WIDTH-1:0] wire_d32_53;
	wire [WIDTH-1:0] wire_d32_54;
	wire [WIDTH-1:0] wire_d32_55;
	wire [WIDTH-1:0] wire_d32_56;
	wire [WIDTH-1:0] wire_d32_57;
	wire [WIDTH-1:0] wire_d32_58;
	wire [WIDTH-1:0] wire_d32_59;
	wire [WIDTH-1:0] wire_d32_60;
	wire [WIDTH-1:0] wire_d32_61;
	wire [WIDTH-1:0] wire_d32_62;
	wire [WIDTH-1:0] wire_d32_63;
	wire [WIDTH-1:0] wire_d32_64;
	wire [WIDTH-1:0] wire_d32_65;
	wire [WIDTH-1:0] wire_d32_66;
	wire [WIDTH-1:0] wire_d32_67;
	wire [WIDTH-1:0] wire_d32_68;
	wire [WIDTH-1:0] wire_d32_69;
	wire [WIDTH-1:0] wire_d32_70;
	wire [WIDTH-1:0] wire_d32_71;
	wire [WIDTH-1:0] wire_d32_72;
	wire [WIDTH-1:0] wire_d32_73;
	wire [WIDTH-1:0] wire_d32_74;
	wire [WIDTH-1:0] wire_d32_75;
	wire [WIDTH-1:0] wire_d32_76;
	wire [WIDTH-1:0] wire_d32_77;
	wire [WIDTH-1:0] wire_d32_78;
	wire [WIDTH-1:0] wire_d33_0;
	wire [WIDTH-1:0] wire_d33_1;
	wire [WIDTH-1:0] wire_d33_2;
	wire [WIDTH-1:0] wire_d33_3;
	wire [WIDTH-1:0] wire_d33_4;
	wire [WIDTH-1:0] wire_d33_5;
	wire [WIDTH-1:0] wire_d33_6;
	wire [WIDTH-1:0] wire_d33_7;
	wire [WIDTH-1:0] wire_d33_8;
	wire [WIDTH-1:0] wire_d33_9;
	wire [WIDTH-1:0] wire_d33_10;
	wire [WIDTH-1:0] wire_d33_11;
	wire [WIDTH-1:0] wire_d33_12;
	wire [WIDTH-1:0] wire_d33_13;
	wire [WIDTH-1:0] wire_d33_14;
	wire [WIDTH-1:0] wire_d33_15;
	wire [WIDTH-1:0] wire_d33_16;
	wire [WIDTH-1:0] wire_d33_17;
	wire [WIDTH-1:0] wire_d33_18;
	wire [WIDTH-1:0] wire_d33_19;
	wire [WIDTH-1:0] wire_d33_20;
	wire [WIDTH-1:0] wire_d33_21;
	wire [WIDTH-1:0] wire_d33_22;
	wire [WIDTH-1:0] wire_d33_23;
	wire [WIDTH-1:0] wire_d33_24;
	wire [WIDTH-1:0] wire_d33_25;
	wire [WIDTH-1:0] wire_d33_26;
	wire [WIDTH-1:0] wire_d33_27;
	wire [WIDTH-1:0] wire_d33_28;
	wire [WIDTH-1:0] wire_d33_29;
	wire [WIDTH-1:0] wire_d33_30;
	wire [WIDTH-1:0] wire_d33_31;
	wire [WIDTH-1:0] wire_d33_32;
	wire [WIDTH-1:0] wire_d33_33;
	wire [WIDTH-1:0] wire_d33_34;
	wire [WIDTH-1:0] wire_d33_35;
	wire [WIDTH-1:0] wire_d33_36;
	wire [WIDTH-1:0] wire_d33_37;
	wire [WIDTH-1:0] wire_d33_38;
	wire [WIDTH-1:0] wire_d33_39;
	wire [WIDTH-1:0] wire_d33_40;
	wire [WIDTH-1:0] wire_d33_41;
	wire [WIDTH-1:0] wire_d33_42;
	wire [WIDTH-1:0] wire_d33_43;
	wire [WIDTH-1:0] wire_d33_44;
	wire [WIDTH-1:0] wire_d33_45;
	wire [WIDTH-1:0] wire_d33_46;
	wire [WIDTH-1:0] wire_d33_47;
	wire [WIDTH-1:0] wire_d33_48;
	wire [WIDTH-1:0] wire_d33_49;
	wire [WIDTH-1:0] wire_d33_50;
	wire [WIDTH-1:0] wire_d33_51;
	wire [WIDTH-1:0] wire_d33_52;
	wire [WIDTH-1:0] wire_d33_53;
	wire [WIDTH-1:0] wire_d33_54;
	wire [WIDTH-1:0] wire_d33_55;
	wire [WIDTH-1:0] wire_d33_56;
	wire [WIDTH-1:0] wire_d33_57;
	wire [WIDTH-1:0] wire_d33_58;
	wire [WIDTH-1:0] wire_d33_59;
	wire [WIDTH-1:0] wire_d33_60;
	wire [WIDTH-1:0] wire_d33_61;
	wire [WIDTH-1:0] wire_d33_62;
	wire [WIDTH-1:0] wire_d33_63;
	wire [WIDTH-1:0] wire_d33_64;
	wire [WIDTH-1:0] wire_d33_65;
	wire [WIDTH-1:0] wire_d33_66;
	wire [WIDTH-1:0] wire_d33_67;
	wire [WIDTH-1:0] wire_d33_68;
	wire [WIDTH-1:0] wire_d33_69;
	wire [WIDTH-1:0] wire_d33_70;
	wire [WIDTH-1:0] wire_d33_71;
	wire [WIDTH-1:0] wire_d33_72;
	wire [WIDTH-1:0] wire_d33_73;
	wire [WIDTH-1:0] wire_d33_74;
	wire [WIDTH-1:0] wire_d33_75;
	wire [WIDTH-1:0] wire_d33_76;
	wire [WIDTH-1:0] wire_d33_77;
	wire [WIDTH-1:0] wire_d33_78;
	wire [WIDTH-1:0] wire_d34_0;
	wire [WIDTH-1:0] wire_d34_1;
	wire [WIDTH-1:0] wire_d34_2;
	wire [WIDTH-1:0] wire_d34_3;
	wire [WIDTH-1:0] wire_d34_4;
	wire [WIDTH-1:0] wire_d34_5;
	wire [WIDTH-1:0] wire_d34_6;
	wire [WIDTH-1:0] wire_d34_7;
	wire [WIDTH-1:0] wire_d34_8;
	wire [WIDTH-1:0] wire_d34_9;
	wire [WIDTH-1:0] wire_d34_10;
	wire [WIDTH-1:0] wire_d34_11;
	wire [WIDTH-1:0] wire_d34_12;
	wire [WIDTH-1:0] wire_d34_13;
	wire [WIDTH-1:0] wire_d34_14;
	wire [WIDTH-1:0] wire_d34_15;
	wire [WIDTH-1:0] wire_d34_16;
	wire [WIDTH-1:0] wire_d34_17;
	wire [WIDTH-1:0] wire_d34_18;
	wire [WIDTH-1:0] wire_d34_19;
	wire [WIDTH-1:0] wire_d34_20;
	wire [WIDTH-1:0] wire_d34_21;
	wire [WIDTH-1:0] wire_d34_22;
	wire [WIDTH-1:0] wire_d34_23;
	wire [WIDTH-1:0] wire_d34_24;
	wire [WIDTH-1:0] wire_d34_25;
	wire [WIDTH-1:0] wire_d34_26;
	wire [WIDTH-1:0] wire_d34_27;
	wire [WIDTH-1:0] wire_d34_28;
	wire [WIDTH-1:0] wire_d34_29;
	wire [WIDTH-1:0] wire_d34_30;
	wire [WIDTH-1:0] wire_d34_31;
	wire [WIDTH-1:0] wire_d34_32;
	wire [WIDTH-1:0] wire_d34_33;
	wire [WIDTH-1:0] wire_d34_34;
	wire [WIDTH-1:0] wire_d34_35;
	wire [WIDTH-1:0] wire_d34_36;
	wire [WIDTH-1:0] wire_d34_37;
	wire [WIDTH-1:0] wire_d34_38;
	wire [WIDTH-1:0] wire_d34_39;
	wire [WIDTH-1:0] wire_d34_40;
	wire [WIDTH-1:0] wire_d34_41;
	wire [WIDTH-1:0] wire_d34_42;
	wire [WIDTH-1:0] wire_d34_43;
	wire [WIDTH-1:0] wire_d34_44;
	wire [WIDTH-1:0] wire_d34_45;
	wire [WIDTH-1:0] wire_d34_46;
	wire [WIDTH-1:0] wire_d34_47;
	wire [WIDTH-1:0] wire_d34_48;
	wire [WIDTH-1:0] wire_d34_49;
	wire [WIDTH-1:0] wire_d34_50;
	wire [WIDTH-1:0] wire_d34_51;
	wire [WIDTH-1:0] wire_d34_52;
	wire [WIDTH-1:0] wire_d34_53;
	wire [WIDTH-1:0] wire_d34_54;
	wire [WIDTH-1:0] wire_d34_55;
	wire [WIDTH-1:0] wire_d34_56;
	wire [WIDTH-1:0] wire_d34_57;
	wire [WIDTH-1:0] wire_d34_58;
	wire [WIDTH-1:0] wire_d34_59;
	wire [WIDTH-1:0] wire_d34_60;
	wire [WIDTH-1:0] wire_d34_61;
	wire [WIDTH-1:0] wire_d34_62;
	wire [WIDTH-1:0] wire_d34_63;
	wire [WIDTH-1:0] wire_d34_64;
	wire [WIDTH-1:0] wire_d34_65;
	wire [WIDTH-1:0] wire_d34_66;
	wire [WIDTH-1:0] wire_d34_67;
	wire [WIDTH-1:0] wire_d34_68;
	wire [WIDTH-1:0] wire_d34_69;
	wire [WIDTH-1:0] wire_d34_70;
	wire [WIDTH-1:0] wire_d34_71;
	wire [WIDTH-1:0] wire_d34_72;
	wire [WIDTH-1:0] wire_d34_73;
	wire [WIDTH-1:0] wire_d34_74;
	wire [WIDTH-1:0] wire_d34_75;
	wire [WIDTH-1:0] wire_d34_76;
	wire [WIDTH-1:0] wire_d34_77;
	wire [WIDTH-1:0] wire_d34_78;
	wire [WIDTH-1:0] wire_d35_0;
	wire [WIDTH-1:0] wire_d35_1;
	wire [WIDTH-1:0] wire_d35_2;
	wire [WIDTH-1:0] wire_d35_3;
	wire [WIDTH-1:0] wire_d35_4;
	wire [WIDTH-1:0] wire_d35_5;
	wire [WIDTH-1:0] wire_d35_6;
	wire [WIDTH-1:0] wire_d35_7;
	wire [WIDTH-1:0] wire_d35_8;
	wire [WIDTH-1:0] wire_d35_9;
	wire [WIDTH-1:0] wire_d35_10;
	wire [WIDTH-1:0] wire_d35_11;
	wire [WIDTH-1:0] wire_d35_12;
	wire [WIDTH-1:0] wire_d35_13;
	wire [WIDTH-1:0] wire_d35_14;
	wire [WIDTH-1:0] wire_d35_15;
	wire [WIDTH-1:0] wire_d35_16;
	wire [WIDTH-1:0] wire_d35_17;
	wire [WIDTH-1:0] wire_d35_18;
	wire [WIDTH-1:0] wire_d35_19;
	wire [WIDTH-1:0] wire_d35_20;
	wire [WIDTH-1:0] wire_d35_21;
	wire [WIDTH-1:0] wire_d35_22;
	wire [WIDTH-1:0] wire_d35_23;
	wire [WIDTH-1:0] wire_d35_24;
	wire [WIDTH-1:0] wire_d35_25;
	wire [WIDTH-1:0] wire_d35_26;
	wire [WIDTH-1:0] wire_d35_27;
	wire [WIDTH-1:0] wire_d35_28;
	wire [WIDTH-1:0] wire_d35_29;
	wire [WIDTH-1:0] wire_d35_30;
	wire [WIDTH-1:0] wire_d35_31;
	wire [WIDTH-1:0] wire_d35_32;
	wire [WIDTH-1:0] wire_d35_33;
	wire [WIDTH-1:0] wire_d35_34;
	wire [WIDTH-1:0] wire_d35_35;
	wire [WIDTH-1:0] wire_d35_36;
	wire [WIDTH-1:0] wire_d35_37;
	wire [WIDTH-1:0] wire_d35_38;
	wire [WIDTH-1:0] wire_d35_39;
	wire [WIDTH-1:0] wire_d35_40;
	wire [WIDTH-1:0] wire_d35_41;
	wire [WIDTH-1:0] wire_d35_42;
	wire [WIDTH-1:0] wire_d35_43;
	wire [WIDTH-1:0] wire_d35_44;
	wire [WIDTH-1:0] wire_d35_45;
	wire [WIDTH-1:0] wire_d35_46;
	wire [WIDTH-1:0] wire_d35_47;
	wire [WIDTH-1:0] wire_d35_48;
	wire [WIDTH-1:0] wire_d35_49;
	wire [WIDTH-1:0] wire_d35_50;
	wire [WIDTH-1:0] wire_d35_51;
	wire [WIDTH-1:0] wire_d35_52;
	wire [WIDTH-1:0] wire_d35_53;
	wire [WIDTH-1:0] wire_d35_54;
	wire [WIDTH-1:0] wire_d35_55;
	wire [WIDTH-1:0] wire_d35_56;
	wire [WIDTH-1:0] wire_d35_57;
	wire [WIDTH-1:0] wire_d35_58;
	wire [WIDTH-1:0] wire_d35_59;
	wire [WIDTH-1:0] wire_d35_60;
	wire [WIDTH-1:0] wire_d35_61;
	wire [WIDTH-1:0] wire_d35_62;
	wire [WIDTH-1:0] wire_d35_63;
	wire [WIDTH-1:0] wire_d35_64;
	wire [WIDTH-1:0] wire_d35_65;
	wire [WIDTH-1:0] wire_d35_66;
	wire [WIDTH-1:0] wire_d35_67;
	wire [WIDTH-1:0] wire_d35_68;
	wire [WIDTH-1:0] wire_d35_69;
	wire [WIDTH-1:0] wire_d35_70;
	wire [WIDTH-1:0] wire_d35_71;
	wire [WIDTH-1:0] wire_d35_72;
	wire [WIDTH-1:0] wire_d35_73;
	wire [WIDTH-1:0] wire_d35_74;
	wire [WIDTH-1:0] wire_d35_75;
	wire [WIDTH-1:0] wire_d35_76;
	wire [WIDTH-1:0] wire_d35_77;
	wire [WIDTH-1:0] wire_d35_78;
	wire [WIDTH-1:0] wire_d36_0;
	wire [WIDTH-1:0] wire_d36_1;
	wire [WIDTH-1:0] wire_d36_2;
	wire [WIDTH-1:0] wire_d36_3;
	wire [WIDTH-1:0] wire_d36_4;
	wire [WIDTH-1:0] wire_d36_5;
	wire [WIDTH-1:0] wire_d36_6;
	wire [WIDTH-1:0] wire_d36_7;
	wire [WIDTH-1:0] wire_d36_8;
	wire [WIDTH-1:0] wire_d36_9;
	wire [WIDTH-1:0] wire_d36_10;
	wire [WIDTH-1:0] wire_d36_11;
	wire [WIDTH-1:0] wire_d36_12;
	wire [WIDTH-1:0] wire_d36_13;
	wire [WIDTH-1:0] wire_d36_14;
	wire [WIDTH-1:0] wire_d36_15;
	wire [WIDTH-1:0] wire_d36_16;
	wire [WIDTH-1:0] wire_d36_17;
	wire [WIDTH-1:0] wire_d36_18;
	wire [WIDTH-1:0] wire_d36_19;
	wire [WIDTH-1:0] wire_d36_20;
	wire [WIDTH-1:0] wire_d36_21;
	wire [WIDTH-1:0] wire_d36_22;
	wire [WIDTH-1:0] wire_d36_23;
	wire [WIDTH-1:0] wire_d36_24;
	wire [WIDTH-1:0] wire_d36_25;
	wire [WIDTH-1:0] wire_d36_26;
	wire [WIDTH-1:0] wire_d36_27;
	wire [WIDTH-1:0] wire_d36_28;
	wire [WIDTH-1:0] wire_d36_29;
	wire [WIDTH-1:0] wire_d36_30;
	wire [WIDTH-1:0] wire_d36_31;
	wire [WIDTH-1:0] wire_d36_32;
	wire [WIDTH-1:0] wire_d36_33;
	wire [WIDTH-1:0] wire_d36_34;
	wire [WIDTH-1:0] wire_d36_35;
	wire [WIDTH-1:0] wire_d36_36;
	wire [WIDTH-1:0] wire_d36_37;
	wire [WIDTH-1:0] wire_d36_38;
	wire [WIDTH-1:0] wire_d36_39;
	wire [WIDTH-1:0] wire_d36_40;
	wire [WIDTH-1:0] wire_d36_41;
	wire [WIDTH-1:0] wire_d36_42;
	wire [WIDTH-1:0] wire_d36_43;
	wire [WIDTH-1:0] wire_d36_44;
	wire [WIDTH-1:0] wire_d36_45;
	wire [WIDTH-1:0] wire_d36_46;
	wire [WIDTH-1:0] wire_d36_47;
	wire [WIDTH-1:0] wire_d36_48;
	wire [WIDTH-1:0] wire_d36_49;
	wire [WIDTH-1:0] wire_d36_50;
	wire [WIDTH-1:0] wire_d36_51;
	wire [WIDTH-1:0] wire_d36_52;
	wire [WIDTH-1:0] wire_d36_53;
	wire [WIDTH-1:0] wire_d36_54;
	wire [WIDTH-1:0] wire_d36_55;
	wire [WIDTH-1:0] wire_d36_56;
	wire [WIDTH-1:0] wire_d36_57;
	wire [WIDTH-1:0] wire_d36_58;
	wire [WIDTH-1:0] wire_d36_59;
	wire [WIDTH-1:0] wire_d36_60;
	wire [WIDTH-1:0] wire_d36_61;
	wire [WIDTH-1:0] wire_d36_62;
	wire [WIDTH-1:0] wire_d36_63;
	wire [WIDTH-1:0] wire_d36_64;
	wire [WIDTH-1:0] wire_d36_65;
	wire [WIDTH-1:0] wire_d36_66;
	wire [WIDTH-1:0] wire_d36_67;
	wire [WIDTH-1:0] wire_d36_68;
	wire [WIDTH-1:0] wire_d36_69;
	wire [WIDTH-1:0] wire_d36_70;
	wire [WIDTH-1:0] wire_d36_71;
	wire [WIDTH-1:0] wire_d36_72;
	wire [WIDTH-1:0] wire_d36_73;
	wire [WIDTH-1:0] wire_d36_74;
	wire [WIDTH-1:0] wire_d36_75;
	wire [WIDTH-1:0] wire_d36_76;
	wire [WIDTH-1:0] wire_d36_77;
	wire [WIDTH-1:0] wire_d36_78;
	wire [WIDTH-1:0] wire_d37_0;
	wire [WIDTH-1:0] wire_d37_1;
	wire [WIDTH-1:0] wire_d37_2;
	wire [WIDTH-1:0] wire_d37_3;
	wire [WIDTH-1:0] wire_d37_4;
	wire [WIDTH-1:0] wire_d37_5;
	wire [WIDTH-1:0] wire_d37_6;
	wire [WIDTH-1:0] wire_d37_7;
	wire [WIDTH-1:0] wire_d37_8;
	wire [WIDTH-1:0] wire_d37_9;
	wire [WIDTH-1:0] wire_d37_10;
	wire [WIDTH-1:0] wire_d37_11;
	wire [WIDTH-1:0] wire_d37_12;
	wire [WIDTH-1:0] wire_d37_13;
	wire [WIDTH-1:0] wire_d37_14;
	wire [WIDTH-1:0] wire_d37_15;
	wire [WIDTH-1:0] wire_d37_16;
	wire [WIDTH-1:0] wire_d37_17;
	wire [WIDTH-1:0] wire_d37_18;
	wire [WIDTH-1:0] wire_d37_19;
	wire [WIDTH-1:0] wire_d37_20;
	wire [WIDTH-1:0] wire_d37_21;
	wire [WIDTH-1:0] wire_d37_22;
	wire [WIDTH-1:0] wire_d37_23;
	wire [WIDTH-1:0] wire_d37_24;
	wire [WIDTH-1:0] wire_d37_25;
	wire [WIDTH-1:0] wire_d37_26;
	wire [WIDTH-1:0] wire_d37_27;
	wire [WIDTH-1:0] wire_d37_28;
	wire [WIDTH-1:0] wire_d37_29;
	wire [WIDTH-1:0] wire_d37_30;
	wire [WIDTH-1:0] wire_d37_31;
	wire [WIDTH-1:0] wire_d37_32;
	wire [WIDTH-1:0] wire_d37_33;
	wire [WIDTH-1:0] wire_d37_34;
	wire [WIDTH-1:0] wire_d37_35;
	wire [WIDTH-1:0] wire_d37_36;
	wire [WIDTH-1:0] wire_d37_37;
	wire [WIDTH-1:0] wire_d37_38;
	wire [WIDTH-1:0] wire_d37_39;
	wire [WIDTH-1:0] wire_d37_40;
	wire [WIDTH-1:0] wire_d37_41;
	wire [WIDTH-1:0] wire_d37_42;
	wire [WIDTH-1:0] wire_d37_43;
	wire [WIDTH-1:0] wire_d37_44;
	wire [WIDTH-1:0] wire_d37_45;
	wire [WIDTH-1:0] wire_d37_46;
	wire [WIDTH-1:0] wire_d37_47;
	wire [WIDTH-1:0] wire_d37_48;
	wire [WIDTH-1:0] wire_d37_49;
	wire [WIDTH-1:0] wire_d37_50;
	wire [WIDTH-1:0] wire_d37_51;
	wire [WIDTH-1:0] wire_d37_52;
	wire [WIDTH-1:0] wire_d37_53;
	wire [WIDTH-1:0] wire_d37_54;
	wire [WIDTH-1:0] wire_d37_55;
	wire [WIDTH-1:0] wire_d37_56;
	wire [WIDTH-1:0] wire_d37_57;
	wire [WIDTH-1:0] wire_d37_58;
	wire [WIDTH-1:0] wire_d37_59;
	wire [WIDTH-1:0] wire_d37_60;
	wire [WIDTH-1:0] wire_d37_61;
	wire [WIDTH-1:0] wire_d37_62;
	wire [WIDTH-1:0] wire_d37_63;
	wire [WIDTH-1:0] wire_d37_64;
	wire [WIDTH-1:0] wire_d37_65;
	wire [WIDTH-1:0] wire_d37_66;
	wire [WIDTH-1:0] wire_d37_67;
	wire [WIDTH-1:0] wire_d37_68;
	wire [WIDTH-1:0] wire_d37_69;
	wire [WIDTH-1:0] wire_d37_70;
	wire [WIDTH-1:0] wire_d37_71;
	wire [WIDTH-1:0] wire_d37_72;
	wire [WIDTH-1:0] wire_d37_73;
	wire [WIDTH-1:0] wire_d37_74;
	wire [WIDTH-1:0] wire_d37_75;
	wire [WIDTH-1:0] wire_d37_76;
	wire [WIDTH-1:0] wire_d37_77;
	wire [WIDTH-1:0] wire_d37_78;
	wire [WIDTH-1:0] wire_d38_0;
	wire [WIDTH-1:0] wire_d38_1;
	wire [WIDTH-1:0] wire_d38_2;
	wire [WIDTH-1:0] wire_d38_3;
	wire [WIDTH-1:0] wire_d38_4;
	wire [WIDTH-1:0] wire_d38_5;
	wire [WIDTH-1:0] wire_d38_6;
	wire [WIDTH-1:0] wire_d38_7;
	wire [WIDTH-1:0] wire_d38_8;
	wire [WIDTH-1:0] wire_d38_9;
	wire [WIDTH-1:0] wire_d38_10;
	wire [WIDTH-1:0] wire_d38_11;
	wire [WIDTH-1:0] wire_d38_12;
	wire [WIDTH-1:0] wire_d38_13;
	wire [WIDTH-1:0] wire_d38_14;
	wire [WIDTH-1:0] wire_d38_15;
	wire [WIDTH-1:0] wire_d38_16;
	wire [WIDTH-1:0] wire_d38_17;
	wire [WIDTH-1:0] wire_d38_18;
	wire [WIDTH-1:0] wire_d38_19;
	wire [WIDTH-1:0] wire_d38_20;
	wire [WIDTH-1:0] wire_d38_21;
	wire [WIDTH-1:0] wire_d38_22;
	wire [WIDTH-1:0] wire_d38_23;
	wire [WIDTH-1:0] wire_d38_24;
	wire [WIDTH-1:0] wire_d38_25;
	wire [WIDTH-1:0] wire_d38_26;
	wire [WIDTH-1:0] wire_d38_27;
	wire [WIDTH-1:0] wire_d38_28;
	wire [WIDTH-1:0] wire_d38_29;
	wire [WIDTH-1:0] wire_d38_30;
	wire [WIDTH-1:0] wire_d38_31;
	wire [WIDTH-1:0] wire_d38_32;
	wire [WIDTH-1:0] wire_d38_33;
	wire [WIDTH-1:0] wire_d38_34;
	wire [WIDTH-1:0] wire_d38_35;
	wire [WIDTH-1:0] wire_d38_36;
	wire [WIDTH-1:0] wire_d38_37;
	wire [WIDTH-1:0] wire_d38_38;
	wire [WIDTH-1:0] wire_d38_39;
	wire [WIDTH-1:0] wire_d38_40;
	wire [WIDTH-1:0] wire_d38_41;
	wire [WIDTH-1:0] wire_d38_42;
	wire [WIDTH-1:0] wire_d38_43;
	wire [WIDTH-1:0] wire_d38_44;
	wire [WIDTH-1:0] wire_d38_45;
	wire [WIDTH-1:0] wire_d38_46;
	wire [WIDTH-1:0] wire_d38_47;
	wire [WIDTH-1:0] wire_d38_48;
	wire [WIDTH-1:0] wire_d38_49;
	wire [WIDTH-1:0] wire_d38_50;
	wire [WIDTH-1:0] wire_d38_51;
	wire [WIDTH-1:0] wire_d38_52;
	wire [WIDTH-1:0] wire_d38_53;
	wire [WIDTH-1:0] wire_d38_54;
	wire [WIDTH-1:0] wire_d38_55;
	wire [WIDTH-1:0] wire_d38_56;
	wire [WIDTH-1:0] wire_d38_57;
	wire [WIDTH-1:0] wire_d38_58;
	wire [WIDTH-1:0] wire_d38_59;
	wire [WIDTH-1:0] wire_d38_60;
	wire [WIDTH-1:0] wire_d38_61;
	wire [WIDTH-1:0] wire_d38_62;
	wire [WIDTH-1:0] wire_d38_63;
	wire [WIDTH-1:0] wire_d38_64;
	wire [WIDTH-1:0] wire_d38_65;
	wire [WIDTH-1:0] wire_d38_66;
	wire [WIDTH-1:0] wire_d38_67;
	wire [WIDTH-1:0] wire_d38_68;
	wire [WIDTH-1:0] wire_d38_69;
	wire [WIDTH-1:0] wire_d38_70;
	wire [WIDTH-1:0] wire_d38_71;
	wire [WIDTH-1:0] wire_d38_72;
	wire [WIDTH-1:0] wire_d38_73;
	wire [WIDTH-1:0] wire_d38_74;
	wire [WIDTH-1:0] wire_d38_75;
	wire [WIDTH-1:0] wire_d38_76;
	wire [WIDTH-1:0] wire_d38_77;
	wire [WIDTH-1:0] wire_d38_78;
	wire [WIDTH-1:0] wire_d39_0;
	wire [WIDTH-1:0] wire_d39_1;
	wire [WIDTH-1:0] wire_d39_2;
	wire [WIDTH-1:0] wire_d39_3;
	wire [WIDTH-1:0] wire_d39_4;
	wire [WIDTH-1:0] wire_d39_5;
	wire [WIDTH-1:0] wire_d39_6;
	wire [WIDTH-1:0] wire_d39_7;
	wire [WIDTH-1:0] wire_d39_8;
	wire [WIDTH-1:0] wire_d39_9;
	wire [WIDTH-1:0] wire_d39_10;
	wire [WIDTH-1:0] wire_d39_11;
	wire [WIDTH-1:0] wire_d39_12;
	wire [WIDTH-1:0] wire_d39_13;
	wire [WIDTH-1:0] wire_d39_14;
	wire [WIDTH-1:0] wire_d39_15;
	wire [WIDTH-1:0] wire_d39_16;
	wire [WIDTH-1:0] wire_d39_17;
	wire [WIDTH-1:0] wire_d39_18;
	wire [WIDTH-1:0] wire_d39_19;
	wire [WIDTH-1:0] wire_d39_20;
	wire [WIDTH-1:0] wire_d39_21;
	wire [WIDTH-1:0] wire_d39_22;
	wire [WIDTH-1:0] wire_d39_23;
	wire [WIDTH-1:0] wire_d39_24;
	wire [WIDTH-1:0] wire_d39_25;
	wire [WIDTH-1:0] wire_d39_26;
	wire [WIDTH-1:0] wire_d39_27;
	wire [WIDTH-1:0] wire_d39_28;
	wire [WIDTH-1:0] wire_d39_29;
	wire [WIDTH-1:0] wire_d39_30;
	wire [WIDTH-1:0] wire_d39_31;
	wire [WIDTH-1:0] wire_d39_32;
	wire [WIDTH-1:0] wire_d39_33;
	wire [WIDTH-1:0] wire_d39_34;
	wire [WIDTH-1:0] wire_d39_35;
	wire [WIDTH-1:0] wire_d39_36;
	wire [WIDTH-1:0] wire_d39_37;
	wire [WIDTH-1:0] wire_d39_38;
	wire [WIDTH-1:0] wire_d39_39;
	wire [WIDTH-1:0] wire_d39_40;
	wire [WIDTH-1:0] wire_d39_41;
	wire [WIDTH-1:0] wire_d39_42;
	wire [WIDTH-1:0] wire_d39_43;
	wire [WIDTH-1:0] wire_d39_44;
	wire [WIDTH-1:0] wire_d39_45;
	wire [WIDTH-1:0] wire_d39_46;
	wire [WIDTH-1:0] wire_d39_47;
	wire [WIDTH-1:0] wire_d39_48;
	wire [WIDTH-1:0] wire_d39_49;
	wire [WIDTH-1:0] wire_d39_50;
	wire [WIDTH-1:0] wire_d39_51;
	wire [WIDTH-1:0] wire_d39_52;
	wire [WIDTH-1:0] wire_d39_53;
	wire [WIDTH-1:0] wire_d39_54;
	wire [WIDTH-1:0] wire_d39_55;
	wire [WIDTH-1:0] wire_d39_56;
	wire [WIDTH-1:0] wire_d39_57;
	wire [WIDTH-1:0] wire_d39_58;
	wire [WIDTH-1:0] wire_d39_59;
	wire [WIDTH-1:0] wire_d39_60;
	wire [WIDTH-1:0] wire_d39_61;
	wire [WIDTH-1:0] wire_d39_62;
	wire [WIDTH-1:0] wire_d39_63;
	wire [WIDTH-1:0] wire_d39_64;
	wire [WIDTH-1:0] wire_d39_65;
	wire [WIDTH-1:0] wire_d39_66;
	wire [WIDTH-1:0] wire_d39_67;
	wire [WIDTH-1:0] wire_d39_68;
	wire [WIDTH-1:0] wire_d39_69;
	wire [WIDTH-1:0] wire_d39_70;
	wire [WIDTH-1:0] wire_d39_71;
	wire [WIDTH-1:0] wire_d39_72;
	wire [WIDTH-1:0] wire_d39_73;
	wire [WIDTH-1:0] wire_d39_74;
	wire [WIDTH-1:0] wire_d39_75;
	wire [WIDTH-1:0] wire_d39_76;
	wire [WIDTH-1:0] wire_d39_77;
	wire [WIDTH-1:0] wire_d39_78;
	wire [WIDTH-1:0] wire_d40_0;
	wire [WIDTH-1:0] wire_d40_1;
	wire [WIDTH-1:0] wire_d40_2;
	wire [WIDTH-1:0] wire_d40_3;
	wire [WIDTH-1:0] wire_d40_4;
	wire [WIDTH-1:0] wire_d40_5;
	wire [WIDTH-1:0] wire_d40_6;
	wire [WIDTH-1:0] wire_d40_7;
	wire [WIDTH-1:0] wire_d40_8;
	wire [WIDTH-1:0] wire_d40_9;
	wire [WIDTH-1:0] wire_d40_10;
	wire [WIDTH-1:0] wire_d40_11;
	wire [WIDTH-1:0] wire_d40_12;
	wire [WIDTH-1:0] wire_d40_13;
	wire [WIDTH-1:0] wire_d40_14;
	wire [WIDTH-1:0] wire_d40_15;
	wire [WIDTH-1:0] wire_d40_16;
	wire [WIDTH-1:0] wire_d40_17;
	wire [WIDTH-1:0] wire_d40_18;
	wire [WIDTH-1:0] wire_d40_19;
	wire [WIDTH-1:0] wire_d40_20;
	wire [WIDTH-1:0] wire_d40_21;
	wire [WIDTH-1:0] wire_d40_22;
	wire [WIDTH-1:0] wire_d40_23;
	wire [WIDTH-1:0] wire_d40_24;
	wire [WIDTH-1:0] wire_d40_25;
	wire [WIDTH-1:0] wire_d40_26;
	wire [WIDTH-1:0] wire_d40_27;
	wire [WIDTH-1:0] wire_d40_28;
	wire [WIDTH-1:0] wire_d40_29;
	wire [WIDTH-1:0] wire_d40_30;
	wire [WIDTH-1:0] wire_d40_31;
	wire [WIDTH-1:0] wire_d40_32;
	wire [WIDTH-1:0] wire_d40_33;
	wire [WIDTH-1:0] wire_d40_34;
	wire [WIDTH-1:0] wire_d40_35;
	wire [WIDTH-1:0] wire_d40_36;
	wire [WIDTH-1:0] wire_d40_37;
	wire [WIDTH-1:0] wire_d40_38;
	wire [WIDTH-1:0] wire_d40_39;
	wire [WIDTH-1:0] wire_d40_40;
	wire [WIDTH-1:0] wire_d40_41;
	wire [WIDTH-1:0] wire_d40_42;
	wire [WIDTH-1:0] wire_d40_43;
	wire [WIDTH-1:0] wire_d40_44;
	wire [WIDTH-1:0] wire_d40_45;
	wire [WIDTH-1:0] wire_d40_46;
	wire [WIDTH-1:0] wire_d40_47;
	wire [WIDTH-1:0] wire_d40_48;
	wire [WIDTH-1:0] wire_d40_49;
	wire [WIDTH-1:0] wire_d40_50;
	wire [WIDTH-1:0] wire_d40_51;
	wire [WIDTH-1:0] wire_d40_52;
	wire [WIDTH-1:0] wire_d40_53;
	wire [WIDTH-1:0] wire_d40_54;
	wire [WIDTH-1:0] wire_d40_55;
	wire [WIDTH-1:0] wire_d40_56;
	wire [WIDTH-1:0] wire_d40_57;
	wire [WIDTH-1:0] wire_d40_58;
	wire [WIDTH-1:0] wire_d40_59;
	wire [WIDTH-1:0] wire_d40_60;
	wire [WIDTH-1:0] wire_d40_61;
	wire [WIDTH-1:0] wire_d40_62;
	wire [WIDTH-1:0] wire_d40_63;
	wire [WIDTH-1:0] wire_d40_64;
	wire [WIDTH-1:0] wire_d40_65;
	wire [WIDTH-1:0] wire_d40_66;
	wire [WIDTH-1:0] wire_d40_67;
	wire [WIDTH-1:0] wire_d40_68;
	wire [WIDTH-1:0] wire_d40_69;
	wire [WIDTH-1:0] wire_d40_70;
	wire [WIDTH-1:0] wire_d40_71;
	wire [WIDTH-1:0] wire_d40_72;
	wire [WIDTH-1:0] wire_d40_73;
	wire [WIDTH-1:0] wire_d40_74;
	wire [WIDTH-1:0] wire_d40_75;
	wire [WIDTH-1:0] wire_d40_76;
	wire [WIDTH-1:0] wire_d40_77;
	wire [WIDTH-1:0] wire_d40_78;
	wire [WIDTH-1:0] wire_d41_0;
	wire [WIDTH-1:0] wire_d41_1;
	wire [WIDTH-1:0] wire_d41_2;
	wire [WIDTH-1:0] wire_d41_3;
	wire [WIDTH-1:0] wire_d41_4;
	wire [WIDTH-1:0] wire_d41_5;
	wire [WIDTH-1:0] wire_d41_6;
	wire [WIDTH-1:0] wire_d41_7;
	wire [WIDTH-1:0] wire_d41_8;
	wire [WIDTH-1:0] wire_d41_9;
	wire [WIDTH-1:0] wire_d41_10;
	wire [WIDTH-1:0] wire_d41_11;
	wire [WIDTH-1:0] wire_d41_12;
	wire [WIDTH-1:0] wire_d41_13;
	wire [WIDTH-1:0] wire_d41_14;
	wire [WIDTH-1:0] wire_d41_15;
	wire [WIDTH-1:0] wire_d41_16;
	wire [WIDTH-1:0] wire_d41_17;
	wire [WIDTH-1:0] wire_d41_18;
	wire [WIDTH-1:0] wire_d41_19;
	wire [WIDTH-1:0] wire_d41_20;
	wire [WIDTH-1:0] wire_d41_21;
	wire [WIDTH-1:0] wire_d41_22;
	wire [WIDTH-1:0] wire_d41_23;
	wire [WIDTH-1:0] wire_d41_24;
	wire [WIDTH-1:0] wire_d41_25;
	wire [WIDTH-1:0] wire_d41_26;
	wire [WIDTH-1:0] wire_d41_27;
	wire [WIDTH-1:0] wire_d41_28;
	wire [WIDTH-1:0] wire_d41_29;
	wire [WIDTH-1:0] wire_d41_30;
	wire [WIDTH-1:0] wire_d41_31;
	wire [WIDTH-1:0] wire_d41_32;
	wire [WIDTH-1:0] wire_d41_33;
	wire [WIDTH-1:0] wire_d41_34;
	wire [WIDTH-1:0] wire_d41_35;
	wire [WIDTH-1:0] wire_d41_36;
	wire [WIDTH-1:0] wire_d41_37;
	wire [WIDTH-1:0] wire_d41_38;
	wire [WIDTH-1:0] wire_d41_39;
	wire [WIDTH-1:0] wire_d41_40;
	wire [WIDTH-1:0] wire_d41_41;
	wire [WIDTH-1:0] wire_d41_42;
	wire [WIDTH-1:0] wire_d41_43;
	wire [WIDTH-1:0] wire_d41_44;
	wire [WIDTH-1:0] wire_d41_45;
	wire [WIDTH-1:0] wire_d41_46;
	wire [WIDTH-1:0] wire_d41_47;
	wire [WIDTH-1:0] wire_d41_48;
	wire [WIDTH-1:0] wire_d41_49;
	wire [WIDTH-1:0] wire_d41_50;
	wire [WIDTH-1:0] wire_d41_51;
	wire [WIDTH-1:0] wire_d41_52;
	wire [WIDTH-1:0] wire_d41_53;
	wire [WIDTH-1:0] wire_d41_54;
	wire [WIDTH-1:0] wire_d41_55;
	wire [WIDTH-1:0] wire_d41_56;
	wire [WIDTH-1:0] wire_d41_57;
	wire [WIDTH-1:0] wire_d41_58;
	wire [WIDTH-1:0] wire_d41_59;
	wire [WIDTH-1:0] wire_d41_60;
	wire [WIDTH-1:0] wire_d41_61;
	wire [WIDTH-1:0] wire_d41_62;
	wire [WIDTH-1:0] wire_d41_63;
	wire [WIDTH-1:0] wire_d41_64;
	wire [WIDTH-1:0] wire_d41_65;
	wire [WIDTH-1:0] wire_d41_66;
	wire [WIDTH-1:0] wire_d41_67;
	wire [WIDTH-1:0] wire_d41_68;
	wire [WIDTH-1:0] wire_d41_69;
	wire [WIDTH-1:0] wire_d41_70;
	wire [WIDTH-1:0] wire_d41_71;
	wire [WIDTH-1:0] wire_d41_72;
	wire [WIDTH-1:0] wire_d41_73;
	wire [WIDTH-1:0] wire_d41_74;
	wire [WIDTH-1:0] wire_d41_75;
	wire [WIDTH-1:0] wire_d41_76;
	wire [WIDTH-1:0] wire_d41_77;
	wire [WIDTH-1:0] wire_d41_78;
	wire [WIDTH-1:0] wire_d42_0;
	wire [WIDTH-1:0] wire_d42_1;
	wire [WIDTH-1:0] wire_d42_2;
	wire [WIDTH-1:0] wire_d42_3;
	wire [WIDTH-1:0] wire_d42_4;
	wire [WIDTH-1:0] wire_d42_5;
	wire [WIDTH-1:0] wire_d42_6;
	wire [WIDTH-1:0] wire_d42_7;
	wire [WIDTH-1:0] wire_d42_8;
	wire [WIDTH-1:0] wire_d42_9;
	wire [WIDTH-1:0] wire_d42_10;
	wire [WIDTH-1:0] wire_d42_11;
	wire [WIDTH-1:0] wire_d42_12;
	wire [WIDTH-1:0] wire_d42_13;
	wire [WIDTH-1:0] wire_d42_14;
	wire [WIDTH-1:0] wire_d42_15;
	wire [WIDTH-1:0] wire_d42_16;
	wire [WIDTH-1:0] wire_d42_17;
	wire [WIDTH-1:0] wire_d42_18;
	wire [WIDTH-1:0] wire_d42_19;
	wire [WIDTH-1:0] wire_d42_20;
	wire [WIDTH-1:0] wire_d42_21;
	wire [WIDTH-1:0] wire_d42_22;
	wire [WIDTH-1:0] wire_d42_23;
	wire [WIDTH-1:0] wire_d42_24;
	wire [WIDTH-1:0] wire_d42_25;
	wire [WIDTH-1:0] wire_d42_26;
	wire [WIDTH-1:0] wire_d42_27;
	wire [WIDTH-1:0] wire_d42_28;
	wire [WIDTH-1:0] wire_d42_29;
	wire [WIDTH-1:0] wire_d42_30;
	wire [WIDTH-1:0] wire_d42_31;
	wire [WIDTH-1:0] wire_d42_32;
	wire [WIDTH-1:0] wire_d42_33;
	wire [WIDTH-1:0] wire_d42_34;
	wire [WIDTH-1:0] wire_d42_35;
	wire [WIDTH-1:0] wire_d42_36;
	wire [WIDTH-1:0] wire_d42_37;
	wire [WIDTH-1:0] wire_d42_38;
	wire [WIDTH-1:0] wire_d42_39;
	wire [WIDTH-1:0] wire_d42_40;
	wire [WIDTH-1:0] wire_d42_41;
	wire [WIDTH-1:0] wire_d42_42;
	wire [WIDTH-1:0] wire_d42_43;
	wire [WIDTH-1:0] wire_d42_44;
	wire [WIDTH-1:0] wire_d42_45;
	wire [WIDTH-1:0] wire_d42_46;
	wire [WIDTH-1:0] wire_d42_47;
	wire [WIDTH-1:0] wire_d42_48;
	wire [WIDTH-1:0] wire_d42_49;
	wire [WIDTH-1:0] wire_d42_50;
	wire [WIDTH-1:0] wire_d42_51;
	wire [WIDTH-1:0] wire_d42_52;
	wire [WIDTH-1:0] wire_d42_53;
	wire [WIDTH-1:0] wire_d42_54;
	wire [WIDTH-1:0] wire_d42_55;
	wire [WIDTH-1:0] wire_d42_56;
	wire [WIDTH-1:0] wire_d42_57;
	wire [WIDTH-1:0] wire_d42_58;
	wire [WIDTH-1:0] wire_d42_59;
	wire [WIDTH-1:0] wire_d42_60;
	wire [WIDTH-1:0] wire_d42_61;
	wire [WIDTH-1:0] wire_d42_62;
	wire [WIDTH-1:0] wire_d42_63;
	wire [WIDTH-1:0] wire_d42_64;
	wire [WIDTH-1:0] wire_d42_65;
	wire [WIDTH-1:0] wire_d42_66;
	wire [WIDTH-1:0] wire_d42_67;
	wire [WIDTH-1:0] wire_d42_68;
	wire [WIDTH-1:0] wire_d42_69;
	wire [WIDTH-1:0] wire_d42_70;
	wire [WIDTH-1:0] wire_d42_71;
	wire [WIDTH-1:0] wire_d42_72;
	wire [WIDTH-1:0] wire_d42_73;
	wire [WIDTH-1:0] wire_d42_74;
	wire [WIDTH-1:0] wire_d42_75;
	wire [WIDTH-1:0] wire_d42_76;
	wire [WIDTH-1:0] wire_d42_77;
	wire [WIDTH-1:0] wire_d42_78;
	wire [WIDTH-1:0] wire_d43_0;
	wire [WIDTH-1:0] wire_d43_1;
	wire [WIDTH-1:0] wire_d43_2;
	wire [WIDTH-1:0] wire_d43_3;
	wire [WIDTH-1:0] wire_d43_4;
	wire [WIDTH-1:0] wire_d43_5;
	wire [WIDTH-1:0] wire_d43_6;
	wire [WIDTH-1:0] wire_d43_7;
	wire [WIDTH-1:0] wire_d43_8;
	wire [WIDTH-1:0] wire_d43_9;
	wire [WIDTH-1:0] wire_d43_10;
	wire [WIDTH-1:0] wire_d43_11;
	wire [WIDTH-1:0] wire_d43_12;
	wire [WIDTH-1:0] wire_d43_13;
	wire [WIDTH-1:0] wire_d43_14;
	wire [WIDTH-1:0] wire_d43_15;
	wire [WIDTH-1:0] wire_d43_16;
	wire [WIDTH-1:0] wire_d43_17;
	wire [WIDTH-1:0] wire_d43_18;
	wire [WIDTH-1:0] wire_d43_19;
	wire [WIDTH-1:0] wire_d43_20;
	wire [WIDTH-1:0] wire_d43_21;
	wire [WIDTH-1:0] wire_d43_22;
	wire [WIDTH-1:0] wire_d43_23;
	wire [WIDTH-1:0] wire_d43_24;
	wire [WIDTH-1:0] wire_d43_25;
	wire [WIDTH-1:0] wire_d43_26;
	wire [WIDTH-1:0] wire_d43_27;
	wire [WIDTH-1:0] wire_d43_28;
	wire [WIDTH-1:0] wire_d43_29;
	wire [WIDTH-1:0] wire_d43_30;
	wire [WIDTH-1:0] wire_d43_31;
	wire [WIDTH-1:0] wire_d43_32;
	wire [WIDTH-1:0] wire_d43_33;
	wire [WIDTH-1:0] wire_d43_34;
	wire [WIDTH-1:0] wire_d43_35;
	wire [WIDTH-1:0] wire_d43_36;
	wire [WIDTH-1:0] wire_d43_37;
	wire [WIDTH-1:0] wire_d43_38;
	wire [WIDTH-1:0] wire_d43_39;
	wire [WIDTH-1:0] wire_d43_40;
	wire [WIDTH-1:0] wire_d43_41;
	wire [WIDTH-1:0] wire_d43_42;
	wire [WIDTH-1:0] wire_d43_43;
	wire [WIDTH-1:0] wire_d43_44;
	wire [WIDTH-1:0] wire_d43_45;
	wire [WIDTH-1:0] wire_d43_46;
	wire [WIDTH-1:0] wire_d43_47;
	wire [WIDTH-1:0] wire_d43_48;
	wire [WIDTH-1:0] wire_d43_49;
	wire [WIDTH-1:0] wire_d43_50;
	wire [WIDTH-1:0] wire_d43_51;
	wire [WIDTH-1:0] wire_d43_52;
	wire [WIDTH-1:0] wire_d43_53;
	wire [WIDTH-1:0] wire_d43_54;
	wire [WIDTH-1:0] wire_d43_55;
	wire [WIDTH-1:0] wire_d43_56;
	wire [WIDTH-1:0] wire_d43_57;
	wire [WIDTH-1:0] wire_d43_58;
	wire [WIDTH-1:0] wire_d43_59;
	wire [WIDTH-1:0] wire_d43_60;
	wire [WIDTH-1:0] wire_d43_61;
	wire [WIDTH-1:0] wire_d43_62;
	wire [WIDTH-1:0] wire_d43_63;
	wire [WIDTH-1:0] wire_d43_64;
	wire [WIDTH-1:0] wire_d43_65;
	wire [WIDTH-1:0] wire_d43_66;
	wire [WIDTH-1:0] wire_d43_67;
	wire [WIDTH-1:0] wire_d43_68;
	wire [WIDTH-1:0] wire_d43_69;
	wire [WIDTH-1:0] wire_d43_70;
	wire [WIDTH-1:0] wire_d43_71;
	wire [WIDTH-1:0] wire_d43_72;
	wire [WIDTH-1:0] wire_d43_73;
	wire [WIDTH-1:0] wire_d43_74;
	wire [WIDTH-1:0] wire_d43_75;
	wire [WIDTH-1:0] wire_d43_76;
	wire [WIDTH-1:0] wire_d43_77;
	wire [WIDTH-1:0] wire_d43_78;
	wire [WIDTH-1:0] wire_d44_0;
	wire [WIDTH-1:0] wire_d44_1;
	wire [WIDTH-1:0] wire_d44_2;
	wire [WIDTH-1:0] wire_d44_3;
	wire [WIDTH-1:0] wire_d44_4;
	wire [WIDTH-1:0] wire_d44_5;
	wire [WIDTH-1:0] wire_d44_6;
	wire [WIDTH-1:0] wire_d44_7;
	wire [WIDTH-1:0] wire_d44_8;
	wire [WIDTH-1:0] wire_d44_9;
	wire [WIDTH-1:0] wire_d44_10;
	wire [WIDTH-1:0] wire_d44_11;
	wire [WIDTH-1:0] wire_d44_12;
	wire [WIDTH-1:0] wire_d44_13;
	wire [WIDTH-1:0] wire_d44_14;
	wire [WIDTH-1:0] wire_d44_15;
	wire [WIDTH-1:0] wire_d44_16;
	wire [WIDTH-1:0] wire_d44_17;
	wire [WIDTH-1:0] wire_d44_18;
	wire [WIDTH-1:0] wire_d44_19;
	wire [WIDTH-1:0] wire_d44_20;
	wire [WIDTH-1:0] wire_d44_21;
	wire [WIDTH-1:0] wire_d44_22;
	wire [WIDTH-1:0] wire_d44_23;
	wire [WIDTH-1:0] wire_d44_24;
	wire [WIDTH-1:0] wire_d44_25;
	wire [WIDTH-1:0] wire_d44_26;
	wire [WIDTH-1:0] wire_d44_27;
	wire [WIDTH-1:0] wire_d44_28;
	wire [WIDTH-1:0] wire_d44_29;
	wire [WIDTH-1:0] wire_d44_30;
	wire [WIDTH-1:0] wire_d44_31;
	wire [WIDTH-1:0] wire_d44_32;
	wire [WIDTH-1:0] wire_d44_33;
	wire [WIDTH-1:0] wire_d44_34;
	wire [WIDTH-1:0] wire_d44_35;
	wire [WIDTH-1:0] wire_d44_36;
	wire [WIDTH-1:0] wire_d44_37;
	wire [WIDTH-1:0] wire_d44_38;
	wire [WIDTH-1:0] wire_d44_39;
	wire [WIDTH-1:0] wire_d44_40;
	wire [WIDTH-1:0] wire_d44_41;
	wire [WIDTH-1:0] wire_d44_42;
	wire [WIDTH-1:0] wire_d44_43;
	wire [WIDTH-1:0] wire_d44_44;
	wire [WIDTH-1:0] wire_d44_45;
	wire [WIDTH-1:0] wire_d44_46;
	wire [WIDTH-1:0] wire_d44_47;
	wire [WIDTH-1:0] wire_d44_48;
	wire [WIDTH-1:0] wire_d44_49;
	wire [WIDTH-1:0] wire_d44_50;
	wire [WIDTH-1:0] wire_d44_51;
	wire [WIDTH-1:0] wire_d44_52;
	wire [WIDTH-1:0] wire_d44_53;
	wire [WIDTH-1:0] wire_d44_54;
	wire [WIDTH-1:0] wire_d44_55;
	wire [WIDTH-1:0] wire_d44_56;
	wire [WIDTH-1:0] wire_d44_57;
	wire [WIDTH-1:0] wire_d44_58;
	wire [WIDTH-1:0] wire_d44_59;
	wire [WIDTH-1:0] wire_d44_60;
	wire [WIDTH-1:0] wire_d44_61;
	wire [WIDTH-1:0] wire_d44_62;
	wire [WIDTH-1:0] wire_d44_63;
	wire [WIDTH-1:0] wire_d44_64;
	wire [WIDTH-1:0] wire_d44_65;
	wire [WIDTH-1:0] wire_d44_66;
	wire [WIDTH-1:0] wire_d44_67;
	wire [WIDTH-1:0] wire_d44_68;
	wire [WIDTH-1:0] wire_d44_69;
	wire [WIDTH-1:0] wire_d44_70;
	wire [WIDTH-1:0] wire_d44_71;
	wire [WIDTH-1:0] wire_d44_72;
	wire [WIDTH-1:0] wire_d44_73;
	wire [WIDTH-1:0] wire_d44_74;
	wire [WIDTH-1:0] wire_d44_75;
	wire [WIDTH-1:0] wire_d44_76;
	wire [WIDTH-1:0] wire_d44_77;
	wire [WIDTH-1:0] wire_d44_78;
	wire [WIDTH-1:0] wire_d45_0;
	wire [WIDTH-1:0] wire_d45_1;
	wire [WIDTH-1:0] wire_d45_2;
	wire [WIDTH-1:0] wire_d45_3;
	wire [WIDTH-1:0] wire_d45_4;
	wire [WIDTH-1:0] wire_d45_5;
	wire [WIDTH-1:0] wire_d45_6;
	wire [WIDTH-1:0] wire_d45_7;
	wire [WIDTH-1:0] wire_d45_8;
	wire [WIDTH-1:0] wire_d45_9;
	wire [WIDTH-1:0] wire_d45_10;
	wire [WIDTH-1:0] wire_d45_11;
	wire [WIDTH-1:0] wire_d45_12;
	wire [WIDTH-1:0] wire_d45_13;
	wire [WIDTH-1:0] wire_d45_14;
	wire [WIDTH-1:0] wire_d45_15;
	wire [WIDTH-1:0] wire_d45_16;
	wire [WIDTH-1:0] wire_d45_17;
	wire [WIDTH-1:0] wire_d45_18;
	wire [WIDTH-1:0] wire_d45_19;
	wire [WIDTH-1:0] wire_d45_20;
	wire [WIDTH-1:0] wire_d45_21;
	wire [WIDTH-1:0] wire_d45_22;
	wire [WIDTH-1:0] wire_d45_23;
	wire [WIDTH-1:0] wire_d45_24;
	wire [WIDTH-1:0] wire_d45_25;
	wire [WIDTH-1:0] wire_d45_26;
	wire [WIDTH-1:0] wire_d45_27;
	wire [WIDTH-1:0] wire_d45_28;
	wire [WIDTH-1:0] wire_d45_29;
	wire [WIDTH-1:0] wire_d45_30;
	wire [WIDTH-1:0] wire_d45_31;
	wire [WIDTH-1:0] wire_d45_32;
	wire [WIDTH-1:0] wire_d45_33;
	wire [WIDTH-1:0] wire_d45_34;
	wire [WIDTH-1:0] wire_d45_35;
	wire [WIDTH-1:0] wire_d45_36;
	wire [WIDTH-1:0] wire_d45_37;
	wire [WIDTH-1:0] wire_d45_38;
	wire [WIDTH-1:0] wire_d45_39;
	wire [WIDTH-1:0] wire_d45_40;
	wire [WIDTH-1:0] wire_d45_41;
	wire [WIDTH-1:0] wire_d45_42;
	wire [WIDTH-1:0] wire_d45_43;
	wire [WIDTH-1:0] wire_d45_44;
	wire [WIDTH-1:0] wire_d45_45;
	wire [WIDTH-1:0] wire_d45_46;
	wire [WIDTH-1:0] wire_d45_47;
	wire [WIDTH-1:0] wire_d45_48;
	wire [WIDTH-1:0] wire_d45_49;
	wire [WIDTH-1:0] wire_d45_50;
	wire [WIDTH-1:0] wire_d45_51;
	wire [WIDTH-1:0] wire_d45_52;
	wire [WIDTH-1:0] wire_d45_53;
	wire [WIDTH-1:0] wire_d45_54;
	wire [WIDTH-1:0] wire_d45_55;
	wire [WIDTH-1:0] wire_d45_56;
	wire [WIDTH-1:0] wire_d45_57;
	wire [WIDTH-1:0] wire_d45_58;
	wire [WIDTH-1:0] wire_d45_59;
	wire [WIDTH-1:0] wire_d45_60;
	wire [WIDTH-1:0] wire_d45_61;
	wire [WIDTH-1:0] wire_d45_62;
	wire [WIDTH-1:0] wire_d45_63;
	wire [WIDTH-1:0] wire_d45_64;
	wire [WIDTH-1:0] wire_d45_65;
	wire [WIDTH-1:0] wire_d45_66;
	wire [WIDTH-1:0] wire_d45_67;
	wire [WIDTH-1:0] wire_d45_68;
	wire [WIDTH-1:0] wire_d45_69;
	wire [WIDTH-1:0] wire_d45_70;
	wire [WIDTH-1:0] wire_d45_71;
	wire [WIDTH-1:0] wire_d45_72;
	wire [WIDTH-1:0] wire_d45_73;
	wire [WIDTH-1:0] wire_d45_74;
	wire [WIDTH-1:0] wire_d45_75;
	wire [WIDTH-1:0] wire_d45_76;
	wire [WIDTH-1:0] wire_d45_77;
	wire [WIDTH-1:0] wire_d45_78;
	wire [WIDTH-1:0] wire_d46_0;
	wire [WIDTH-1:0] wire_d46_1;
	wire [WIDTH-1:0] wire_d46_2;
	wire [WIDTH-1:0] wire_d46_3;
	wire [WIDTH-1:0] wire_d46_4;
	wire [WIDTH-1:0] wire_d46_5;
	wire [WIDTH-1:0] wire_d46_6;
	wire [WIDTH-1:0] wire_d46_7;
	wire [WIDTH-1:0] wire_d46_8;
	wire [WIDTH-1:0] wire_d46_9;
	wire [WIDTH-1:0] wire_d46_10;
	wire [WIDTH-1:0] wire_d46_11;
	wire [WIDTH-1:0] wire_d46_12;
	wire [WIDTH-1:0] wire_d46_13;
	wire [WIDTH-1:0] wire_d46_14;
	wire [WIDTH-1:0] wire_d46_15;
	wire [WIDTH-1:0] wire_d46_16;
	wire [WIDTH-1:0] wire_d46_17;
	wire [WIDTH-1:0] wire_d46_18;
	wire [WIDTH-1:0] wire_d46_19;
	wire [WIDTH-1:0] wire_d46_20;
	wire [WIDTH-1:0] wire_d46_21;
	wire [WIDTH-1:0] wire_d46_22;
	wire [WIDTH-1:0] wire_d46_23;
	wire [WIDTH-1:0] wire_d46_24;
	wire [WIDTH-1:0] wire_d46_25;
	wire [WIDTH-1:0] wire_d46_26;
	wire [WIDTH-1:0] wire_d46_27;
	wire [WIDTH-1:0] wire_d46_28;
	wire [WIDTH-1:0] wire_d46_29;
	wire [WIDTH-1:0] wire_d46_30;
	wire [WIDTH-1:0] wire_d46_31;
	wire [WIDTH-1:0] wire_d46_32;
	wire [WIDTH-1:0] wire_d46_33;
	wire [WIDTH-1:0] wire_d46_34;
	wire [WIDTH-1:0] wire_d46_35;
	wire [WIDTH-1:0] wire_d46_36;
	wire [WIDTH-1:0] wire_d46_37;
	wire [WIDTH-1:0] wire_d46_38;
	wire [WIDTH-1:0] wire_d46_39;
	wire [WIDTH-1:0] wire_d46_40;
	wire [WIDTH-1:0] wire_d46_41;
	wire [WIDTH-1:0] wire_d46_42;
	wire [WIDTH-1:0] wire_d46_43;
	wire [WIDTH-1:0] wire_d46_44;
	wire [WIDTH-1:0] wire_d46_45;
	wire [WIDTH-1:0] wire_d46_46;
	wire [WIDTH-1:0] wire_d46_47;
	wire [WIDTH-1:0] wire_d46_48;
	wire [WIDTH-1:0] wire_d46_49;
	wire [WIDTH-1:0] wire_d46_50;
	wire [WIDTH-1:0] wire_d46_51;
	wire [WIDTH-1:0] wire_d46_52;
	wire [WIDTH-1:0] wire_d46_53;
	wire [WIDTH-1:0] wire_d46_54;
	wire [WIDTH-1:0] wire_d46_55;
	wire [WIDTH-1:0] wire_d46_56;
	wire [WIDTH-1:0] wire_d46_57;
	wire [WIDTH-1:0] wire_d46_58;
	wire [WIDTH-1:0] wire_d46_59;
	wire [WIDTH-1:0] wire_d46_60;
	wire [WIDTH-1:0] wire_d46_61;
	wire [WIDTH-1:0] wire_d46_62;
	wire [WIDTH-1:0] wire_d46_63;
	wire [WIDTH-1:0] wire_d46_64;
	wire [WIDTH-1:0] wire_d46_65;
	wire [WIDTH-1:0] wire_d46_66;
	wire [WIDTH-1:0] wire_d46_67;
	wire [WIDTH-1:0] wire_d46_68;
	wire [WIDTH-1:0] wire_d46_69;
	wire [WIDTH-1:0] wire_d46_70;
	wire [WIDTH-1:0] wire_d46_71;
	wire [WIDTH-1:0] wire_d46_72;
	wire [WIDTH-1:0] wire_d46_73;
	wire [WIDTH-1:0] wire_d46_74;
	wire [WIDTH-1:0] wire_d46_75;
	wire [WIDTH-1:0] wire_d46_76;
	wire [WIDTH-1:0] wire_d46_77;
	wire [WIDTH-1:0] wire_d46_78;
	wire [WIDTH-1:0] wire_d47_0;
	wire [WIDTH-1:0] wire_d47_1;
	wire [WIDTH-1:0] wire_d47_2;
	wire [WIDTH-1:0] wire_d47_3;
	wire [WIDTH-1:0] wire_d47_4;
	wire [WIDTH-1:0] wire_d47_5;
	wire [WIDTH-1:0] wire_d47_6;
	wire [WIDTH-1:0] wire_d47_7;
	wire [WIDTH-1:0] wire_d47_8;
	wire [WIDTH-1:0] wire_d47_9;
	wire [WIDTH-1:0] wire_d47_10;
	wire [WIDTH-1:0] wire_d47_11;
	wire [WIDTH-1:0] wire_d47_12;
	wire [WIDTH-1:0] wire_d47_13;
	wire [WIDTH-1:0] wire_d47_14;
	wire [WIDTH-1:0] wire_d47_15;
	wire [WIDTH-1:0] wire_d47_16;
	wire [WIDTH-1:0] wire_d47_17;
	wire [WIDTH-1:0] wire_d47_18;
	wire [WIDTH-1:0] wire_d47_19;
	wire [WIDTH-1:0] wire_d47_20;
	wire [WIDTH-1:0] wire_d47_21;
	wire [WIDTH-1:0] wire_d47_22;
	wire [WIDTH-1:0] wire_d47_23;
	wire [WIDTH-1:0] wire_d47_24;
	wire [WIDTH-1:0] wire_d47_25;
	wire [WIDTH-1:0] wire_d47_26;
	wire [WIDTH-1:0] wire_d47_27;
	wire [WIDTH-1:0] wire_d47_28;
	wire [WIDTH-1:0] wire_d47_29;
	wire [WIDTH-1:0] wire_d47_30;
	wire [WIDTH-1:0] wire_d47_31;
	wire [WIDTH-1:0] wire_d47_32;
	wire [WIDTH-1:0] wire_d47_33;
	wire [WIDTH-1:0] wire_d47_34;
	wire [WIDTH-1:0] wire_d47_35;
	wire [WIDTH-1:0] wire_d47_36;
	wire [WIDTH-1:0] wire_d47_37;
	wire [WIDTH-1:0] wire_d47_38;
	wire [WIDTH-1:0] wire_d47_39;
	wire [WIDTH-1:0] wire_d47_40;
	wire [WIDTH-1:0] wire_d47_41;
	wire [WIDTH-1:0] wire_d47_42;
	wire [WIDTH-1:0] wire_d47_43;
	wire [WIDTH-1:0] wire_d47_44;
	wire [WIDTH-1:0] wire_d47_45;
	wire [WIDTH-1:0] wire_d47_46;
	wire [WIDTH-1:0] wire_d47_47;
	wire [WIDTH-1:0] wire_d47_48;
	wire [WIDTH-1:0] wire_d47_49;
	wire [WIDTH-1:0] wire_d47_50;
	wire [WIDTH-1:0] wire_d47_51;
	wire [WIDTH-1:0] wire_d47_52;
	wire [WIDTH-1:0] wire_d47_53;
	wire [WIDTH-1:0] wire_d47_54;
	wire [WIDTH-1:0] wire_d47_55;
	wire [WIDTH-1:0] wire_d47_56;
	wire [WIDTH-1:0] wire_d47_57;
	wire [WIDTH-1:0] wire_d47_58;
	wire [WIDTH-1:0] wire_d47_59;
	wire [WIDTH-1:0] wire_d47_60;
	wire [WIDTH-1:0] wire_d47_61;
	wire [WIDTH-1:0] wire_d47_62;
	wire [WIDTH-1:0] wire_d47_63;
	wire [WIDTH-1:0] wire_d47_64;
	wire [WIDTH-1:0] wire_d47_65;
	wire [WIDTH-1:0] wire_d47_66;
	wire [WIDTH-1:0] wire_d47_67;
	wire [WIDTH-1:0] wire_d47_68;
	wire [WIDTH-1:0] wire_d47_69;
	wire [WIDTH-1:0] wire_d47_70;
	wire [WIDTH-1:0] wire_d47_71;
	wire [WIDTH-1:0] wire_d47_72;
	wire [WIDTH-1:0] wire_d47_73;
	wire [WIDTH-1:0] wire_d47_74;
	wire [WIDTH-1:0] wire_d47_75;
	wire [WIDTH-1:0] wire_d47_76;
	wire [WIDTH-1:0] wire_d47_77;
	wire [WIDTH-1:0] wire_d47_78;
	wire [WIDTH-1:0] wire_d48_0;
	wire [WIDTH-1:0] wire_d48_1;
	wire [WIDTH-1:0] wire_d48_2;
	wire [WIDTH-1:0] wire_d48_3;
	wire [WIDTH-1:0] wire_d48_4;
	wire [WIDTH-1:0] wire_d48_5;
	wire [WIDTH-1:0] wire_d48_6;
	wire [WIDTH-1:0] wire_d48_7;
	wire [WIDTH-1:0] wire_d48_8;
	wire [WIDTH-1:0] wire_d48_9;
	wire [WIDTH-1:0] wire_d48_10;
	wire [WIDTH-1:0] wire_d48_11;
	wire [WIDTH-1:0] wire_d48_12;
	wire [WIDTH-1:0] wire_d48_13;
	wire [WIDTH-1:0] wire_d48_14;
	wire [WIDTH-1:0] wire_d48_15;
	wire [WIDTH-1:0] wire_d48_16;
	wire [WIDTH-1:0] wire_d48_17;
	wire [WIDTH-1:0] wire_d48_18;
	wire [WIDTH-1:0] wire_d48_19;
	wire [WIDTH-1:0] wire_d48_20;
	wire [WIDTH-1:0] wire_d48_21;
	wire [WIDTH-1:0] wire_d48_22;
	wire [WIDTH-1:0] wire_d48_23;
	wire [WIDTH-1:0] wire_d48_24;
	wire [WIDTH-1:0] wire_d48_25;
	wire [WIDTH-1:0] wire_d48_26;
	wire [WIDTH-1:0] wire_d48_27;
	wire [WIDTH-1:0] wire_d48_28;
	wire [WIDTH-1:0] wire_d48_29;
	wire [WIDTH-1:0] wire_d48_30;
	wire [WIDTH-1:0] wire_d48_31;
	wire [WIDTH-1:0] wire_d48_32;
	wire [WIDTH-1:0] wire_d48_33;
	wire [WIDTH-1:0] wire_d48_34;
	wire [WIDTH-1:0] wire_d48_35;
	wire [WIDTH-1:0] wire_d48_36;
	wire [WIDTH-1:0] wire_d48_37;
	wire [WIDTH-1:0] wire_d48_38;
	wire [WIDTH-1:0] wire_d48_39;
	wire [WIDTH-1:0] wire_d48_40;
	wire [WIDTH-1:0] wire_d48_41;
	wire [WIDTH-1:0] wire_d48_42;
	wire [WIDTH-1:0] wire_d48_43;
	wire [WIDTH-1:0] wire_d48_44;
	wire [WIDTH-1:0] wire_d48_45;
	wire [WIDTH-1:0] wire_d48_46;
	wire [WIDTH-1:0] wire_d48_47;
	wire [WIDTH-1:0] wire_d48_48;
	wire [WIDTH-1:0] wire_d48_49;
	wire [WIDTH-1:0] wire_d48_50;
	wire [WIDTH-1:0] wire_d48_51;
	wire [WIDTH-1:0] wire_d48_52;
	wire [WIDTH-1:0] wire_d48_53;
	wire [WIDTH-1:0] wire_d48_54;
	wire [WIDTH-1:0] wire_d48_55;
	wire [WIDTH-1:0] wire_d48_56;
	wire [WIDTH-1:0] wire_d48_57;
	wire [WIDTH-1:0] wire_d48_58;
	wire [WIDTH-1:0] wire_d48_59;
	wire [WIDTH-1:0] wire_d48_60;
	wire [WIDTH-1:0] wire_d48_61;
	wire [WIDTH-1:0] wire_d48_62;
	wire [WIDTH-1:0] wire_d48_63;
	wire [WIDTH-1:0] wire_d48_64;
	wire [WIDTH-1:0] wire_d48_65;
	wire [WIDTH-1:0] wire_d48_66;
	wire [WIDTH-1:0] wire_d48_67;
	wire [WIDTH-1:0] wire_d48_68;
	wire [WIDTH-1:0] wire_d48_69;
	wire [WIDTH-1:0] wire_d48_70;
	wire [WIDTH-1:0] wire_d48_71;
	wire [WIDTH-1:0] wire_d48_72;
	wire [WIDTH-1:0] wire_d48_73;
	wire [WIDTH-1:0] wire_d48_74;
	wire [WIDTH-1:0] wire_d48_75;
	wire [WIDTH-1:0] wire_d48_76;
	wire [WIDTH-1:0] wire_d48_77;
	wire [WIDTH-1:0] wire_d48_78;
	wire [WIDTH-1:0] wire_d49_0;
	wire [WIDTH-1:0] wire_d49_1;
	wire [WIDTH-1:0] wire_d49_2;
	wire [WIDTH-1:0] wire_d49_3;
	wire [WIDTH-1:0] wire_d49_4;
	wire [WIDTH-1:0] wire_d49_5;
	wire [WIDTH-1:0] wire_d49_6;
	wire [WIDTH-1:0] wire_d49_7;
	wire [WIDTH-1:0] wire_d49_8;
	wire [WIDTH-1:0] wire_d49_9;
	wire [WIDTH-1:0] wire_d49_10;
	wire [WIDTH-1:0] wire_d49_11;
	wire [WIDTH-1:0] wire_d49_12;
	wire [WIDTH-1:0] wire_d49_13;
	wire [WIDTH-1:0] wire_d49_14;
	wire [WIDTH-1:0] wire_d49_15;
	wire [WIDTH-1:0] wire_d49_16;
	wire [WIDTH-1:0] wire_d49_17;
	wire [WIDTH-1:0] wire_d49_18;
	wire [WIDTH-1:0] wire_d49_19;
	wire [WIDTH-1:0] wire_d49_20;
	wire [WIDTH-1:0] wire_d49_21;
	wire [WIDTH-1:0] wire_d49_22;
	wire [WIDTH-1:0] wire_d49_23;
	wire [WIDTH-1:0] wire_d49_24;
	wire [WIDTH-1:0] wire_d49_25;
	wire [WIDTH-1:0] wire_d49_26;
	wire [WIDTH-1:0] wire_d49_27;
	wire [WIDTH-1:0] wire_d49_28;
	wire [WIDTH-1:0] wire_d49_29;
	wire [WIDTH-1:0] wire_d49_30;
	wire [WIDTH-1:0] wire_d49_31;
	wire [WIDTH-1:0] wire_d49_32;
	wire [WIDTH-1:0] wire_d49_33;
	wire [WIDTH-1:0] wire_d49_34;
	wire [WIDTH-1:0] wire_d49_35;
	wire [WIDTH-1:0] wire_d49_36;
	wire [WIDTH-1:0] wire_d49_37;
	wire [WIDTH-1:0] wire_d49_38;
	wire [WIDTH-1:0] wire_d49_39;
	wire [WIDTH-1:0] wire_d49_40;
	wire [WIDTH-1:0] wire_d49_41;
	wire [WIDTH-1:0] wire_d49_42;
	wire [WIDTH-1:0] wire_d49_43;
	wire [WIDTH-1:0] wire_d49_44;
	wire [WIDTH-1:0] wire_d49_45;
	wire [WIDTH-1:0] wire_d49_46;
	wire [WIDTH-1:0] wire_d49_47;
	wire [WIDTH-1:0] wire_d49_48;
	wire [WIDTH-1:0] wire_d49_49;
	wire [WIDTH-1:0] wire_d49_50;
	wire [WIDTH-1:0] wire_d49_51;
	wire [WIDTH-1:0] wire_d49_52;
	wire [WIDTH-1:0] wire_d49_53;
	wire [WIDTH-1:0] wire_d49_54;
	wire [WIDTH-1:0] wire_d49_55;
	wire [WIDTH-1:0] wire_d49_56;
	wire [WIDTH-1:0] wire_d49_57;
	wire [WIDTH-1:0] wire_d49_58;
	wire [WIDTH-1:0] wire_d49_59;
	wire [WIDTH-1:0] wire_d49_60;
	wire [WIDTH-1:0] wire_d49_61;
	wire [WIDTH-1:0] wire_d49_62;
	wire [WIDTH-1:0] wire_d49_63;
	wire [WIDTH-1:0] wire_d49_64;
	wire [WIDTH-1:0] wire_d49_65;
	wire [WIDTH-1:0] wire_d49_66;
	wire [WIDTH-1:0] wire_d49_67;
	wire [WIDTH-1:0] wire_d49_68;
	wire [WIDTH-1:0] wire_d49_69;
	wire [WIDTH-1:0] wire_d49_70;
	wire [WIDTH-1:0] wire_d49_71;
	wire [WIDTH-1:0] wire_d49_72;
	wire [WIDTH-1:0] wire_d49_73;
	wire [WIDTH-1:0] wire_d49_74;
	wire [WIDTH-1:0] wire_d49_75;
	wire [WIDTH-1:0] wire_d49_76;
	wire [WIDTH-1:0] wire_d49_77;
	wire [WIDTH-1:0] wire_d49_78;
	wire [WIDTH-1:0] wire_d50_0;
	wire [WIDTH-1:0] wire_d50_1;
	wire [WIDTH-1:0] wire_d50_2;
	wire [WIDTH-1:0] wire_d50_3;
	wire [WIDTH-1:0] wire_d50_4;
	wire [WIDTH-1:0] wire_d50_5;
	wire [WIDTH-1:0] wire_d50_6;
	wire [WIDTH-1:0] wire_d50_7;
	wire [WIDTH-1:0] wire_d50_8;
	wire [WIDTH-1:0] wire_d50_9;
	wire [WIDTH-1:0] wire_d50_10;
	wire [WIDTH-1:0] wire_d50_11;
	wire [WIDTH-1:0] wire_d50_12;
	wire [WIDTH-1:0] wire_d50_13;
	wire [WIDTH-1:0] wire_d50_14;
	wire [WIDTH-1:0] wire_d50_15;
	wire [WIDTH-1:0] wire_d50_16;
	wire [WIDTH-1:0] wire_d50_17;
	wire [WIDTH-1:0] wire_d50_18;
	wire [WIDTH-1:0] wire_d50_19;
	wire [WIDTH-1:0] wire_d50_20;
	wire [WIDTH-1:0] wire_d50_21;
	wire [WIDTH-1:0] wire_d50_22;
	wire [WIDTH-1:0] wire_d50_23;
	wire [WIDTH-1:0] wire_d50_24;
	wire [WIDTH-1:0] wire_d50_25;
	wire [WIDTH-1:0] wire_d50_26;
	wire [WIDTH-1:0] wire_d50_27;
	wire [WIDTH-1:0] wire_d50_28;
	wire [WIDTH-1:0] wire_d50_29;
	wire [WIDTH-1:0] wire_d50_30;
	wire [WIDTH-1:0] wire_d50_31;
	wire [WIDTH-1:0] wire_d50_32;
	wire [WIDTH-1:0] wire_d50_33;
	wire [WIDTH-1:0] wire_d50_34;
	wire [WIDTH-1:0] wire_d50_35;
	wire [WIDTH-1:0] wire_d50_36;
	wire [WIDTH-1:0] wire_d50_37;
	wire [WIDTH-1:0] wire_d50_38;
	wire [WIDTH-1:0] wire_d50_39;
	wire [WIDTH-1:0] wire_d50_40;
	wire [WIDTH-1:0] wire_d50_41;
	wire [WIDTH-1:0] wire_d50_42;
	wire [WIDTH-1:0] wire_d50_43;
	wire [WIDTH-1:0] wire_d50_44;
	wire [WIDTH-1:0] wire_d50_45;
	wire [WIDTH-1:0] wire_d50_46;
	wire [WIDTH-1:0] wire_d50_47;
	wire [WIDTH-1:0] wire_d50_48;
	wire [WIDTH-1:0] wire_d50_49;
	wire [WIDTH-1:0] wire_d50_50;
	wire [WIDTH-1:0] wire_d50_51;
	wire [WIDTH-1:0] wire_d50_52;
	wire [WIDTH-1:0] wire_d50_53;
	wire [WIDTH-1:0] wire_d50_54;
	wire [WIDTH-1:0] wire_d50_55;
	wire [WIDTH-1:0] wire_d50_56;
	wire [WIDTH-1:0] wire_d50_57;
	wire [WIDTH-1:0] wire_d50_58;
	wire [WIDTH-1:0] wire_d50_59;
	wire [WIDTH-1:0] wire_d50_60;
	wire [WIDTH-1:0] wire_d50_61;
	wire [WIDTH-1:0] wire_d50_62;
	wire [WIDTH-1:0] wire_d50_63;
	wire [WIDTH-1:0] wire_d50_64;
	wire [WIDTH-1:0] wire_d50_65;
	wire [WIDTH-1:0] wire_d50_66;
	wire [WIDTH-1:0] wire_d50_67;
	wire [WIDTH-1:0] wire_d50_68;
	wire [WIDTH-1:0] wire_d50_69;
	wire [WIDTH-1:0] wire_d50_70;
	wire [WIDTH-1:0] wire_d50_71;
	wire [WIDTH-1:0] wire_d50_72;
	wire [WIDTH-1:0] wire_d50_73;
	wire [WIDTH-1:0] wire_d50_74;
	wire [WIDTH-1:0] wire_d50_75;
	wire [WIDTH-1:0] wire_d50_76;
	wire [WIDTH-1:0] wire_d50_77;
	wire [WIDTH-1:0] wire_d50_78;
	wire [WIDTH-1:0] wire_d51_0;
	wire [WIDTH-1:0] wire_d51_1;
	wire [WIDTH-1:0] wire_d51_2;
	wire [WIDTH-1:0] wire_d51_3;
	wire [WIDTH-1:0] wire_d51_4;
	wire [WIDTH-1:0] wire_d51_5;
	wire [WIDTH-1:0] wire_d51_6;
	wire [WIDTH-1:0] wire_d51_7;
	wire [WIDTH-1:0] wire_d51_8;
	wire [WIDTH-1:0] wire_d51_9;
	wire [WIDTH-1:0] wire_d51_10;
	wire [WIDTH-1:0] wire_d51_11;
	wire [WIDTH-1:0] wire_d51_12;
	wire [WIDTH-1:0] wire_d51_13;
	wire [WIDTH-1:0] wire_d51_14;
	wire [WIDTH-1:0] wire_d51_15;
	wire [WIDTH-1:0] wire_d51_16;
	wire [WIDTH-1:0] wire_d51_17;
	wire [WIDTH-1:0] wire_d51_18;
	wire [WIDTH-1:0] wire_d51_19;
	wire [WIDTH-1:0] wire_d51_20;
	wire [WIDTH-1:0] wire_d51_21;
	wire [WIDTH-1:0] wire_d51_22;
	wire [WIDTH-1:0] wire_d51_23;
	wire [WIDTH-1:0] wire_d51_24;
	wire [WIDTH-1:0] wire_d51_25;
	wire [WIDTH-1:0] wire_d51_26;
	wire [WIDTH-1:0] wire_d51_27;
	wire [WIDTH-1:0] wire_d51_28;
	wire [WIDTH-1:0] wire_d51_29;
	wire [WIDTH-1:0] wire_d51_30;
	wire [WIDTH-1:0] wire_d51_31;
	wire [WIDTH-1:0] wire_d51_32;
	wire [WIDTH-1:0] wire_d51_33;
	wire [WIDTH-1:0] wire_d51_34;
	wire [WIDTH-1:0] wire_d51_35;
	wire [WIDTH-1:0] wire_d51_36;
	wire [WIDTH-1:0] wire_d51_37;
	wire [WIDTH-1:0] wire_d51_38;
	wire [WIDTH-1:0] wire_d51_39;
	wire [WIDTH-1:0] wire_d51_40;
	wire [WIDTH-1:0] wire_d51_41;
	wire [WIDTH-1:0] wire_d51_42;
	wire [WIDTH-1:0] wire_d51_43;
	wire [WIDTH-1:0] wire_d51_44;
	wire [WIDTH-1:0] wire_d51_45;
	wire [WIDTH-1:0] wire_d51_46;
	wire [WIDTH-1:0] wire_d51_47;
	wire [WIDTH-1:0] wire_d51_48;
	wire [WIDTH-1:0] wire_d51_49;
	wire [WIDTH-1:0] wire_d51_50;
	wire [WIDTH-1:0] wire_d51_51;
	wire [WIDTH-1:0] wire_d51_52;
	wire [WIDTH-1:0] wire_d51_53;
	wire [WIDTH-1:0] wire_d51_54;
	wire [WIDTH-1:0] wire_d51_55;
	wire [WIDTH-1:0] wire_d51_56;
	wire [WIDTH-1:0] wire_d51_57;
	wire [WIDTH-1:0] wire_d51_58;
	wire [WIDTH-1:0] wire_d51_59;
	wire [WIDTH-1:0] wire_d51_60;
	wire [WIDTH-1:0] wire_d51_61;
	wire [WIDTH-1:0] wire_d51_62;
	wire [WIDTH-1:0] wire_d51_63;
	wire [WIDTH-1:0] wire_d51_64;
	wire [WIDTH-1:0] wire_d51_65;
	wire [WIDTH-1:0] wire_d51_66;
	wire [WIDTH-1:0] wire_d51_67;
	wire [WIDTH-1:0] wire_d51_68;
	wire [WIDTH-1:0] wire_d51_69;
	wire [WIDTH-1:0] wire_d51_70;
	wire [WIDTH-1:0] wire_d51_71;
	wire [WIDTH-1:0] wire_d51_72;
	wire [WIDTH-1:0] wire_d51_73;
	wire [WIDTH-1:0] wire_d51_74;
	wire [WIDTH-1:0] wire_d51_75;
	wire [WIDTH-1:0] wire_d51_76;
	wire [WIDTH-1:0] wire_d51_77;
	wire [WIDTH-1:0] wire_d51_78;
	wire [WIDTH-1:0] wire_d52_0;
	wire [WIDTH-1:0] wire_d52_1;
	wire [WIDTH-1:0] wire_d52_2;
	wire [WIDTH-1:0] wire_d52_3;
	wire [WIDTH-1:0] wire_d52_4;
	wire [WIDTH-1:0] wire_d52_5;
	wire [WIDTH-1:0] wire_d52_6;
	wire [WIDTH-1:0] wire_d52_7;
	wire [WIDTH-1:0] wire_d52_8;
	wire [WIDTH-1:0] wire_d52_9;
	wire [WIDTH-1:0] wire_d52_10;
	wire [WIDTH-1:0] wire_d52_11;
	wire [WIDTH-1:0] wire_d52_12;
	wire [WIDTH-1:0] wire_d52_13;
	wire [WIDTH-1:0] wire_d52_14;
	wire [WIDTH-1:0] wire_d52_15;
	wire [WIDTH-1:0] wire_d52_16;
	wire [WIDTH-1:0] wire_d52_17;
	wire [WIDTH-1:0] wire_d52_18;
	wire [WIDTH-1:0] wire_d52_19;
	wire [WIDTH-1:0] wire_d52_20;
	wire [WIDTH-1:0] wire_d52_21;
	wire [WIDTH-1:0] wire_d52_22;
	wire [WIDTH-1:0] wire_d52_23;
	wire [WIDTH-1:0] wire_d52_24;
	wire [WIDTH-1:0] wire_d52_25;
	wire [WIDTH-1:0] wire_d52_26;
	wire [WIDTH-1:0] wire_d52_27;
	wire [WIDTH-1:0] wire_d52_28;
	wire [WIDTH-1:0] wire_d52_29;
	wire [WIDTH-1:0] wire_d52_30;
	wire [WIDTH-1:0] wire_d52_31;
	wire [WIDTH-1:0] wire_d52_32;
	wire [WIDTH-1:0] wire_d52_33;
	wire [WIDTH-1:0] wire_d52_34;
	wire [WIDTH-1:0] wire_d52_35;
	wire [WIDTH-1:0] wire_d52_36;
	wire [WIDTH-1:0] wire_d52_37;
	wire [WIDTH-1:0] wire_d52_38;
	wire [WIDTH-1:0] wire_d52_39;
	wire [WIDTH-1:0] wire_d52_40;
	wire [WIDTH-1:0] wire_d52_41;
	wire [WIDTH-1:0] wire_d52_42;
	wire [WIDTH-1:0] wire_d52_43;
	wire [WIDTH-1:0] wire_d52_44;
	wire [WIDTH-1:0] wire_d52_45;
	wire [WIDTH-1:0] wire_d52_46;
	wire [WIDTH-1:0] wire_d52_47;
	wire [WIDTH-1:0] wire_d52_48;
	wire [WIDTH-1:0] wire_d52_49;
	wire [WIDTH-1:0] wire_d52_50;
	wire [WIDTH-1:0] wire_d52_51;
	wire [WIDTH-1:0] wire_d52_52;
	wire [WIDTH-1:0] wire_d52_53;
	wire [WIDTH-1:0] wire_d52_54;
	wire [WIDTH-1:0] wire_d52_55;
	wire [WIDTH-1:0] wire_d52_56;
	wire [WIDTH-1:0] wire_d52_57;
	wire [WIDTH-1:0] wire_d52_58;
	wire [WIDTH-1:0] wire_d52_59;
	wire [WIDTH-1:0] wire_d52_60;
	wire [WIDTH-1:0] wire_d52_61;
	wire [WIDTH-1:0] wire_d52_62;
	wire [WIDTH-1:0] wire_d52_63;
	wire [WIDTH-1:0] wire_d52_64;
	wire [WIDTH-1:0] wire_d52_65;
	wire [WIDTH-1:0] wire_d52_66;
	wire [WIDTH-1:0] wire_d52_67;
	wire [WIDTH-1:0] wire_d52_68;
	wire [WIDTH-1:0] wire_d52_69;
	wire [WIDTH-1:0] wire_d52_70;
	wire [WIDTH-1:0] wire_d52_71;
	wire [WIDTH-1:0] wire_d52_72;
	wire [WIDTH-1:0] wire_d52_73;
	wire [WIDTH-1:0] wire_d52_74;
	wire [WIDTH-1:0] wire_d52_75;
	wire [WIDTH-1:0] wire_d52_76;
	wire [WIDTH-1:0] wire_d52_77;
	wire [WIDTH-1:0] wire_d52_78;
	wire [WIDTH-1:0] wire_d53_0;
	wire [WIDTH-1:0] wire_d53_1;
	wire [WIDTH-1:0] wire_d53_2;
	wire [WIDTH-1:0] wire_d53_3;
	wire [WIDTH-1:0] wire_d53_4;
	wire [WIDTH-1:0] wire_d53_5;
	wire [WIDTH-1:0] wire_d53_6;
	wire [WIDTH-1:0] wire_d53_7;
	wire [WIDTH-1:0] wire_d53_8;
	wire [WIDTH-1:0] wire_d53_9;
	wire [WIDTH-1:0] wire_d53_10;
	wire [WIDTH-1:0] wire_d53_11;
	wire [WIDTH-1:0] wire_d53_12;
	wire [WIDTH-1:0] wire_d53_13;
	wire [WIDTH-1:0] wire_d53_14;
	wire [WIDTH-1:0] wire_d53_15;
	wire [WIDTH-1:0] wire_d53_16;
	wire [WIDTH-1:0] wire_d53_17;
	wire [WIDTH-1:0] wire_d53_18;
	wire [WIDTH-1:0] wire_d53_19;
	wire [WIDTH-1:0] wire_d53_20;
	wire [WIDTH-1:0] wire_d53_21;
	wire [WIDTH-1:0] wire_d53_22;
	wire [WIDTH-1:0] wire_d53_23;
	wire [WIDTH-1:0] wire_d53_24;
	wire [WIDTH-1:0] wire_d53_25;
	wire [WIDTH-1:0] wire_d53_26;
	wire [WIDTH-1:0] wire_d53_27;
	wire [WIDTH-1:0] wire_d53_28;
	wire [WIDTH-1:0] wire_d53_29;
	wire [WIDTH-1:0] wire_d53_30;
	wire [WIDTH-1:0] wire_d53_31;
	wire [WIDTH-1:0] wire_d53_32;
	wire [WIDTH-1:0] wire_d53_33;
	wire [WIDTH-1:0] wire_d53_34;
	wire [WIDTH-1:0] wire_d53_35;
	wire [WIDTH-1:0] wire_d53_36;
	wire [WIDTH-1:0] wire_d53_37;
	wire [WIDTH-1:0] wire_d53_38;
	wire [WIDTH-1:0] wire_d53_39;
	wire [WIDTH-1:0] wire_d53_40;
	wire [WIDTH-1:0] wire_d53_41;
	wire [WIDTH-1:0] wire_d53_42;
	wire [WIDTH-1:0] wire_d53_43;
	wire [WIDTH-1:0] wire_d53_44;
	wire [WIDTH-1:0] wire_d53_45;
	wire [WIDTH-1:0] wire_d53_46;
	wire [WIDTH-1:0] wire_d53_47;
	wire [WIDTH-1:0] wire_d53_48;
	wire [WIDTH-1:0] wire_d53_49;
	wire [WIDTH-1:0] wire_d53_50;
	wire [WIDTH-1:0] wire_d53_51;
	wire [WIDTH-1:0] wire_d53_52;
	wire [WIDTH-1:0] wire_d53_53;
	wire [WIDTH-1:0] wire_d53_54;
	wire [WIDTH-1:0] wire_d53_55;
	wire [WIDTH-1:0] wire_d53_56;
	wire [WIDTH-1:0] wire_d53_57;
	wire [WIDTH-1:0] wire_d53_58;
	wire [WIDTH-1:0] wire_d53_59;
	wire [WIDTH-1:0] wire_d53_60;
	wire [WIDTH-1:0] wire_d53_61;
	wire [WIDTH-1:0] wire_d53_62;
	wire [WIDTH-1:0] wire_d53_63;
	wire [WIDTH-1:0] wire_d53_64;
	wire [WIDTH-1:0] wire_d53_65;
	wire [WIDTH-1:0] wire_d53_66;
	wire [WIDTH-1:0] wire_d53_67;
	wire [WIDTH-1:0] wire_d53_68;
	wire [WIDTH-1:0] wire_d53_69;
	wire [WIDTH-1:0] wire_d53_70;
	wire [WIDTH-1:0] wire_d53_71;
	wire [WIDTH-1:0] wire_d53_72;
	wire [WIDTH-1:0] wire_d53_73;
	wire [WIDTH-1:0] wire_d53_74;
	wire [WIDTH-1:0] wire_d53_75;
	wire [WIDTH-1:0] wire_d53_76;
	wire [WIDTH-1:0] wire_d53_77;
	wire [WIDTH-1:0] wire_d53_78;
	wire [WIDTH-1:0] wire_d54_0;
	wire [WIDTH-1:0] wire_d54_1;
	wire [WIDTH-1:0] wire_d54_2;
	wire [WIDTH-1:0] wire_d54_3;
	wire [WIDTH-1:0] wire_d54_4;
	wire [WIDTH-1:0] wire_d54_5;
	wire [WIDTH-1:0] wire_d54_6;
	wire [WIDTH-1:0] wire_d54_7;
	wire [WIDTH-1:0] wire_d54_8;
	wire [WIDTH-1:0] wire_d54_9;
	wire [WIDTH-1:0] wire_d54_10;
	wire [WIDTH-1:0] wire_d54_11;
	wire [WIDTH-1:0] wire_d54_12;
	wire [WIDTH-1:0] wire_d54_13;
	wire [WIDTH-1:0] wire_d54_14;
	wire [WIDTH-1:0] wire_d54_15;
	wire [WIDTH-1:0] wire_d54_16;
	wire [WIDTH-1:0] wire_d54_17;
	wire [WIDTH-1:0] wire_d54_18;
	wire [WIDTH-1:0] wire_d54_19;
	wire [WIDTH-1:0] wire_d54_20;
	wire [WIDTH-1:0] wire_d54_21;
	wire [WIDTH-1:0] wire_d54_22;
	wire [WIDTH-1:0] wire_d54_23;
	wire [WIDTH-1:0] wire_d54_24;
	wire [WIDTH-1:0] wire_d54_25;
	wire [WIDTH-1:0] wire_d54_26;
	wire [WIDTH-1:0] wire_d54_27;
	wire [WIDTH-1:0] wire_d54_28;
	wire [WIDTH-1:0] wire_d54_29;
	wire [WIDTH-1:0] wire_d54_30;
	wire [WIDTH-1:0] wire_d54_31;
	wire [WIDTH-1:0] wire_d54_32;
	wire [WIDTH-1:0] wire_d54_33;
	wire [WIDTH-1:0] wire_d54_34;
	wire [WIDTH-1:0] wire_d54_35;
	wire [WIDTH-1:0] wire_d54_36;
	wire [WIDTH-1:0] wire_d54_37;
	wire [WIDTH-1:0] wire_d54_38;
	wire [WIDTH-1:0] wire_d54_39;
	wire [WIDTH-1:0] wire_d54_40;
	wire [WIDTH-1:0] wire_d54_41;
	wire [WIDTH-1:0] wire_d54_42;
	wire [WIDTH-1:0] wire_d54_43;
	wire [WIDTH-1:0] wire_d54_44;
	wire [WIDTH-1:0] wire_d54_45;
	wire [WIDTH-1:0] wire_d54_46;
	wire [WIDTH-1:0] wire_d54_47;
	wire [WIDTH-1:0] wire_d54_48;
	wire [WIDTH-1:0] wire_d54_49;
	wire [WIDTH-1:0] wire_d54_50;
	wire [WIDTH-1:0] wire_d54_51;
	wire [WIDTH-1:0] wire_d54_52;
	wire [WIDTH-1:0] wire_d54_53;
	wire [WIDTH-1:0] wire_d54_54;
	wire [WIDTH-1:0] wire_d54_55;
	wire [WIDTH-1:0] wire_d54_56;
	wire [WIDTH-1:0] wire_d54_57;
	wire [WIDTH-1:0] wire_d54_58;
	wire [WIDTH-1:0] wire_d54_59;
	wire [WIDTH-1:0] wire_d54_60;
	wire [WIDTH-1:0] wire_d54_61;
	wire [WIDTH-1:0] wire_d54_62;
	wire [WIDTH-1:0] wire_d54_63;
	wire [WIDTH-1:0] wire_d54_64;
	wire [WIDTH-1:0] wire_d54_65;
	wire [WIDTH-1:0] wire_d54_66;
	wire [WIDTH-1:0] wire_d54_67;
	wire [WIDTH-1:0] wire_d54_68;
	wire [WIDTH-1:0] wire_d54_69;
	wire [WIDTH-1:0] wire_d54_70;
	wire [WIDTH-1:0] wire_d54_71;
	wire [WIDTH-1:0] wire_d54_72;
	wire [WIDTH-1:0] wire_d54_73;
	wire [WIDTH-1:0] wire_d54_74;
	wire [WIDTH-1:0] wire_d54_75;
	wire [WIDTH-1:0] wire_d54_76;
	wire [WIDTH-1:0] wire_d54_77;
	wire [WIDTH-1:0] wire_d54_78;
	wire [WIDTH-1:0] wire_d55_0;
	wire [WIDTH-1:0] wire_d55_1;
	wire [WIDTH-1:0] wire_d55_2;
	wire [WIDTH-1:0] wire_d55_3;
	wire [WIDTH-1:0] wire_d55_4;
	wire [WIDTH-1:0] wire_d55_5;
	wire [WIDTH-1:0] wire_d55_6;
	wire [WIDTH-1:0] wire_d55_7;
	wire [WIDTH-1:0] wire_d55_8;
	wire [WIDTH-1:0] wire_d55_9;
	wire [WIDTH-1:0] wire_d55_10;
	wire [WIDTH-1:0] wire_d55_11;
	wire [WIDTH-1:0] wire_d55_12;
	wire [WIDTH-1:0] wire_d55_13;
	wire [WIDTH-1:0] wire_d55_14;
	wire [WIDTH-1:0] wire_d55_15;
	wire [WIDTH-1:0] wire_d55_16;
	wire [WIDTH-1:0] wire_d55_17;
	wire [WIDTH-1:0] wire_d55_18;
	wire [WIDTH-1:0] wire_d55_19;
	wire [WIDTH-1:0] wire_d55_20;
	wire [WIDTH-1:0] wire_d55_21;
	wire [WIDTH-1:0] wire_d55_22;
	wire [WIDTH-1:0] wire_d55_23;
	wire [WIDTH-1:0] wire_d55_24;
	wire [WIDTH-1:0] wire_d55_25;
	wire [WIDTH-1:0] wire_d55_26;
	wire [WIDTH-1:0] wire_d55_27;
	wire [WIDTH-1:0] wire_d55_28;
	wire [WIDTH-1:0] wire_d55_29;
	wire [WIDTH-1:0] wire_d55_30;
	wire [WIDTH-1:0] wire_d55_31;
	wire [WIDTH-1:0] wire_d55_32;
	wire [WIDTH-1:0] wire_d55_33;
	wire [WIDTH-1:0] wire_d55_34;
	wire [WIDTH-1:0] wire_d55_35;
	wire [WIDTH-1:0] wire_d55_36;
	wire [WIDTH-1:0] wire_d55_37;
	wire [WIDTH-1:0] wire_d55_38;
	wire [WIDTH-1:0] wire_d55_39;
	wire [WIDTH-1:0] wire_d55_40;
	wire [WIDTH-1:0] wire_d55_41;
	wire [WIDTH-1:0] wire_d55_42;
	wire [WIDTH-1:0] wire_d55_43;
	wire [WIDTH-1:0] wire_d55_44;
	wire [WIDTH-1:0] wire_d55_45;
	wire [WIDTH-1:0] wire_d55_46;
	wire [WIDTH-1:0] wire_d55_47;
	wire [WIDTH-1:0] wire_d55_48;
	wire [WIDTH-1:0] wire_d55_49;
	wire [WIDTH-1:0] wire_d55_50;
	wire [WIDTH-1:0] wire_d55_51;
	wire [WIDTH-1:0] wire_d55_52;
	wire [WIDTH-1:0] wire_d55_53;
	wire [WIDTH-1:0] wire_d55_54;
	wire [WIDTH-1:0] wire_d55_55;
	wire [WIDTH-1:0] wire_d55_56;
	wire [WIDTH-1:0] wire_d55_57;
	wire [WIDTH-1:0] wire_d55_58;
	wire [WIDTH-1:0] wire_d55_59;
	wire [WIDTH-1:0] wire_d55_60;
	wire [WIDTH-1:0] wire_d55_61;
	wire [WIDTH-1:0] wire_d55_62;
	wire [WIDTH-1:0] wire_d55_63;
	wire [WIDTH-1:0] wire_d55_64;
	wire [WIDTH-1:0] wire_d55_65;
	wire [WIDTH-1:0] wire_d55_66;
	wire [WIDTH-1:0] wire_d55_67;
	wire [WIDTH-1:0] wire_d55_68;
	wire [WIDTH-1:0] wire_d55_69;
	wire [WIDTH-1:0] wire_d55_70;
	wire [WIDTH-1:0] wire_d55_71;
	wire [WIDTH-1:0] wire_d55_72;
	wire [WIDTH-1:0] wire_d55_73;
	wire [WIDTH-1:0] wire_d55_74;
	wire [WIDTH-1:0] wire_d55_75;
	wire [WIDTH-1:0] wire_d55_76;
	wire [WIDTH-1:0] wire_d55_77;
	wire [WIDTH-1:0] wire_d55_78;
	wire [WIDTH-1:0] wire_d56_0;
	wire [WIDTH-1:0] wire_d56_1;
	wire [WIDTH-1:0] wire_d56_2;
	wire [WIDTH-1:0] wire_d56_3;
	wire [WIDTH-1:0] wire_d56_4;
	wire [WIDTH-1:0] wire_d56_5;
	wire [WIDTH-1:0] wire_d56_6;
	wire [WIDTH-1:0] wire_d56_7;
	wire [WIDTH-1:0] wire_d56_8;
	wire [WIDTH-1:0] wire_d56_9;
	wire [WIDTH-1:0] wire_d56_10;
	wire [WIDTH-1:0] wire_d56_11;
	wire [WIDTH-1:0] wire_d56_12;
	wire [WIDTH-1:0] wire_d56_13;
	wire [WIDTH-1:0] wire_d56_14;
	wire [WIDTH-1:0] wire_d56_15;
	wire [WIDTH-1:0] wire_d56_16;
	wire [WIDTH-1:0] wire_d56_17;
	wire [WIDTH-1:0] wire_d56_18;
	wire [WIDTH-1:0] wire_d56_19;
	wire [WIDTH-1:0] wire_d56_20;
	wire [WIDTH-1:0] wire_d56_21;
	wire [WIDTH-1:0] wire_d56_22;
	wire [WIDTH-1:0] wire_d56_23;
	wire [WIDTH-1:0] wire_d56_24;
	wire [WIDTH-1:0] wire_d56_25;
	wire [WIDTH-1:0] wire_d56_26;
	wire [WIDTH-1:0] wire_d56_27;
	wire [WIDTH-1:0] wire_d56_28;
	wire [WIDTH-1:0] wire_d56_29;
	wire [WIDTH-1:0] wire_d56_30;
	wire [WIDTH-1:0] wire_d56_31;
	wire [WIDTH-1:0] wire_d56_32;
	wire [WIDTH-1:0] wire_d56_33;
	wire [WIDTH-1:0] wire_d56_34;
	wire [WIDTH-1:0] wire_d56_35;
	wire [WIDTH-1:0] wire_d56_36;
	wire [WIDTH-1:0] wire_d56_37;
	wire [WIDTH-1:0] wire_d56_38;
	wire [WIDTH-1:0] wire_d56_39;
	wire [WIDTH-1:0] wire_d56_40;
	wire [WIDTH-1:0] wire_d56_41;
	wire [WIDTH-1:0] wire_d56_42;
	wire [WIDTH-1:0] wire_d56_43;
	wire [WIDTH-1:0] wire_d56_44;
	wire [WIDTH-1:0] wire_d56_45;
	wire [WIDTH-1:0] wire_d56_46;
	wire [WIDTH-1:0] wire_d56_47;
	wire [WIDTH-1:0] wire_d56_48;
	wire [WIDTH-1:0] wire_d56_49;
	wire [WIDTH-1:0] wire_d56_50;
	wire [WIDTH-1:0] wire_d56_51;
	wire [WIDTH-1:0] wire_d56_52;
	wire [WIDTH-1:0] wire_d56_53;
	wire [WIDTH-1:0] wire_d56_54;
	wire [WIDTH-1:0] wire_d56_55;
	wire [WIDTH-1:0] wire_d56_56;
	wire [WIDTH-1:0] wire_d56_57;
	wire [WIDTH-1:0] wire_d56_58;
	wire [WIDTH-1:0] wire_d56_59;
	wire [WIDTH-1:0] wire_d56_60;
	wire [WIDTH-1:0] wire_d56_61;
	wire [WIDTH-1:0] wire_d56_62;
	wire [WIDTH-1:0] wire_d56_63;
	wire [WIDTH-1:0] wire_d56_64;
	wire [WIDTH-1:0] wire_d56_65;
	wire [WIDTH-1:0] wire_d56_66;
	wire [WIDTH-1:0] wire_d56_67;
	wire [WIDTH-1:0] wire_d56_68;
	wire [WIDTH-1:0] wire_d56_69;
	wire [WIDTH-1:0] wire_d56_70;
	wire [WIDTH-1:0] wire_d56_71;
	wire [WIDTH-1:0] wire_d56_72;
	wire [WIDTH-1:0] wire_d56_73;
	wire [WIDTH-1:0] wire_d56_74;
	wire [WIDTH-1:0] wire_d56_75;
	wire [WIDTH-1:0] wire_d56_76;
	wire [WIDTH-1:0] wire_d56_77;
	wire [WIDTH-1:0] wire_d56_78;
	wire [WIDTH-1:0] wire_d57_0;
	wire [WIDTH-1:0] wire_d57_1;
	wire [WIDTH-1:0] wire_d57_2;
	wire [WIDTH-1:0] wire_d57_3;
	wire [WIDTH-1:0] wire_d57_4;
	wire [WIDTH-1:0] wire_d57_5;
	wire [WIDTH-1:0] wire_d57_6;
	wire [WIDTH-1:0] wire_d57_7;
	wire [WIDTH-1:0] wire_d57_8;
	wire [WIDTH-1:0] wire_d57_9;
	wire [WIDTH-1:0] wire_d57_10;
	wire [WIDTH-1:0] wire_d57_11;
	wire [WIDTH-1:0] wire_d57_12;
	wire [WIDTH-1:0] wire_d57_13;
	wire [WIDTH-1:0] wire_d57_14;
	wire [WIDTH-1:0] wire_d57_15;
	wire [WIDTH-1:0] wire_d57_16;
	wire [WIDTH-1:0] wire_d57_17;
	wire [WIDTH-1:0] wire_d57_18;
	wire [WIDTH-1:0] wire_d57_19;
	wire [WIDTH-1:0] wire_d57_20;
	wire [WIDTH-1:0] wire_d57_21;
	wire [WIDTH-1:0] wire_d57_22;
	wire [WIDTH-1:0] wire_d57_23;
	wire [WIDTH-1:0] wire_d57_24;
	wire [WIDTH-1:0] wire_d57_25;
	wire [WIDTH-1:0] wire_d57_26;
	wire [WIDTH-1:0] wire_d57_27;
	wire [WIDTH-1:0] wire_d57_28;
	wire [WIDTH-1:0] wire_d57_29;
	wire [WIDTH-1:0] wire_d57_30;
	wire [WIDTH-1:0] wire_d57_31;
	wire [WIDTH-1:0] wire_d57_32;
	wire [WIDTH-1:0] wire_d57_33;
	wire [WIDTH-1:0] wire_d57_34;
	wire [WIDTH-1:0] wire_d57_35;
	wire [WIDTH-1:0] wire_d57_36;
	wire [WIDTH-1:0] wire_d57_37;
	wire [WIDTH-1:0] wire_d57_38;
	wire [WIDTH-1:0] wire_d57_39;
	wire [WIDTH-1:0] wire_d57_40;
	wire [WIDTH-1:0] wire_d57_41;
	wire [WIDTH-1:0] wire_d57_42;
	wire [WIDTH-1:0] wire_d57_43;
	wire [WIDTH-1:0] wire_d57_44;
	wire [WIDTH-1:0] wire_d57_45;
	wire [WIDTH-1:0] wire_d57_46;
	wire [WIDTH-1:0] wire_d57_47;
	wire [WIDTH-1:0] wire_d57_48;
	wire [WIDTH-1:0] wire_d57_49;
	wire [WIDTH-1:0] wire_d57_50;
	wire [WIDTH-1:0] wire_d57_51;
	wire [WIDTH-1:0] wire_d57_52;
	wire [WIDTH-1:0] wire_d57_53;
	wire [WIDTH-1:0] wire_d57_54;
	wire [WIDTH-1:0] wire_d57_55;
	wire [WIDTH-1:0] wire_d57_56;
	wire [WIDTH-1:0] wire_d57_57;
	wire [WIDTH-1:0] wire_d57_58;
	wire [WIDTH-1:0] wire_d57_59;
	wire [WIDTH-1:0] wire_d57_60;
	wire [WIDTH-1:0] wire_d57_61;
	wire [WIDTH-1:0] wire_d57_62;
	wire [WIDTH-1:0] wire_d57_63;
	wire [WIDTH-1:0] wire_d57_64;
	wire [WIDTH-1:0] wire_d57_65;
	wire [WIDTH-1:0] wire_d57_66;
	wire [WIDTH-1:0] wire_d57_67;
	wire [WIDTH-1:0] wire_d57_68;
	wire [WIDTH-1:0] wire_d57_69;
	wire [WIDTH-1:0] wire_d57_70;
	wire [WIDTH-1:0] wire_d57_71;
	wire [WIDTH-1:0] wire_d57_72;
	wire [WIDTH-1:0] wire_d57_73;
	wire [WIDTH-1:0] wire_d57_74;
	wire [WIDTH-1:0] wire_d57_75;
	wire [WIDTH-1:0] wire_d57_76;
	wire [WIDTH-1:0] wire_d57_77;
	wire [WIDTH-1:0] wire_d57_78;
	wire [WIDTH-1:0] wire_d58_0;
	wire [WIDTH-1:0] wire_d58_1;
	wire [WIDTH-1:0] wire_d58_2;
	wire [WIDTH-1:0] wire_d58_3;
	wire [WIDTH-1:0] wire_d58_4;
	wire [WIDTH-1:0] wire_d58_5;
	wire [WIDTH-1:0] wire_d58_6;
	wire [WIDTH-1:0] wire_d58_7;
	wire [WIDTH-1:0] wire_d58_8;
	wire [WIDTH-1:0] wire_d58_9;
	wire [WIDTH-1:0] wire_d58_10;
	wire [WIDTH-1:0] wire_d58_11;
	wire [WIDTH-1:0] wire_d58_12;
	wire [WIDTH-1:0] wire_d58_13;
	wire [WIDTH-1:0] wire_d58_14;
	wire [WIDTH-1:0] wire_d58_15;
	wire [WIDTH-1:0] wire_d58_16;
	wire [WIDTH-1:0] wire_d58_17;
	wire [WIDTH-1:0] wire_d58_18;
	wire [WIDTH-1:0] wire_d58_19;
	wire [WIDTH-1:0] wire_d58_20;
	wire [WIDTH-1:0] wire_d58_21;
	wire [WIDTH-1:0] wire_d58_22;
	wire [WIDTH-1:0] wire_d58_23;
	wire [WIDTH-1:0] wire_d58_24;
	wire [WIDTH-1:0] wire_d58_25;
	wire [WIDTH-1:0] wire_d58_26;
	wire [WIDTH-1:0] wire_d58_27;
	wire [WIDTH-1:0] wire_d58_28;
	wire [WIDTH-1:0] wire_d58_29;
	wire [WIDTH-1:0] wire_d58_30;
	wire [WIDTH-1:0] wire_d58_31;
	wire [WIDTH-1:0] wire_d58_32;
	wire [WIDTH-1:0] wire_d58_33;
	wire [WIDTH-1:0] wire_d58_34;
	wire [WIDTH-1:0] wire_d58_35;
	wire [WIDTH-1:0] wire_d58_36;
	wire [WIDTH-1:0] wire_d58_37;
	wire [WIDTH-1:0] wire_d58_38;
	wire [WIDTH-1:0] wire_d58_39;
	wire [WIDTH-1:0] wire_d58_40;
	wire [WIDTH-1:0] wire_d58_41;
	wire [WIDTH-1:0] wire_d58_42;
	wire [WIDTH-1:0] wire_d58_43;
	wire [WIDTH-1:0] wire_d58_44;
	wire [WIDTH-1:0] wire_d58_45;
	wire [WIDTH-1:0] wire_d58_46;
	wire [WIDTH-1:0] wire_d58_47;
	wire [WIDTH-1:0] wire_d58_48;
	wire [WIDTH-1:0] wire_d58_49;
	wire [WIDTH-1:0] wire_d58_50;
	wire [WIDTH-1:0] wire_d58_51;
	wire [WIDTH-1:0] wire_d58_52;
	wire [WIDTH-1:0] wire_d58_53;
	wire [WIDTH-1:0] wire_d58_54;
	wire [WIDTH-1:0] wire_d58_55;
	wire [WIDTH-1:0] wire_d58_56;
	wire [WIDTH-1:0] wire_d58_57;
	wire [WIDTH-1:0] wire_d58_58;
	wire [WIDTH-1:0] wire_d58_59;
	wire [WIDTH-1:0] wire_d58_60;
	wire [WIDTH-1:0] wire_d58_61;
	wire [WIDTH-1:0] wire_d58_62;
	wire [WIDTH-1:0] wire_d58_63;
	wire [WIDTH-1:0] wire_d58_64;
	wire [WIDTH-1:0] wire_d58_65;
	wire [WIDTH-1:0] wire_d58_66;
	wire [WIDTH-1:0] wire_d58_67;
	wire [WIDTH-1:0] wire_d58_68;
	wire [WIDTH-1:0] wire_d58_69;
	wire [WIDTH-1:0] wire_d58_70;
	wire [WIDTH-1:0] wire_d58_71;
	wire [WIDTH-1:0] wire_d58_72;
	wire [WIDTH-1:0] wire_d58_73;
	wire [WIDTH-1:0] wire_d58_74;
	wire [WIDTH-1:0] wire_d58_75;
	wire [WIDTH-1:0] wire_d58_76;
	wire [WIDTH-1:0] wire_d58_77;
	wire [WIDTH-1:0] wire_d58_78;
	wire [WIDTH-1:0] wire_d59_0;
	wire [WIDTH-1:0] wire_d59_1;
	wire [WIDTH-1:0] wire_d59_2;
	wire [WIDTH-1:0] wire_d59_3;
	wire [WIDTH-1:0] wire_d59_4;
	wire [WIDTH-1:0] wire_d59_5;
	wire [WIDTH-1:0] wire_d59_6;
	wire [WIDTH-1:0] wire_d59_7;
	wire [WIDTH-1:0] wire_d59_8;
	wire [WIDTH-1:0] wire_d59_9;
	wire [WIDTH-1:0] wire_d59_10;
	wire [WIDTH-1:0] wire_d59_11;
	wire [WIDTH-1:0] wire_d59_12;
	wire [WIDTH-1:0] wire_d59_13;
	wire [WIDTH-1:0] wire_d59_14;
	wire [WIDTH-1:0] wire_d59_15;
	wire [WIDTH-1:0] wire_d59_16;
	wire [WIDTH-1:0] wire_d59_17;
	wire [WIDTH-1:0] wire_d59_18;
	wire [WIDTH-1:0] wire_d59_19;
	wire [WIDTH-1:0] wire_d59_20;
	wire [WIDTH-1:0] wire_d59_21;
	wire [WIDTH-1:0] wire_d59_22;
	wire [WIDTH-1:0] wire_d59_23;
	wire [WIDTH-1:0] wire_d59_24;
	wire [WIDTH-1:0] wire_d59_25;
	wire [WIDTH-1:0] wire_d59_26;
	wire [WIDTH-1:0] wire_d59_27;
	wire [WIDTH-1:0] wire_d59_28;
	wire [WIDTH-1:0] wire_d59_29;
	wire [WIDTH-1:0] wire_d59_30;
	wire [WIDTH-1:0] wire_d59_31;
	wire [WIDTH-1:0] wire_d59_32;
	wire [WIDTH-1:0] wire_d59_33;
	wire [WIDTH-1:0] wire_d59_34;
	wire [WIDTH-1:0] wire_d59_35;
	wire [WIDTH-1:0] wire_d59_36;
	wire [WIDTH-1:0] wire_d59_37;
	wire [WIDTH-1:0] wire_d59_38;
	wire [WIDTH-1:0] wire_d59_39;
	wire [WIDTH-1:0] wire_d59_40;
	wire [WIDTH-1:0] wire_d59_41;
	wire [WIDTH-1:0] wire_d59_42;
	wire [WIDTH-1:0] wire_d59_43;
	wire [WIDTH-1:0] wire_d59_44;
	wire [WIDTH-1:0] wire_d59_45;
	wire [WIDTH-1:0] wire_d59_46;
	wire [WIDTH-1:0] wire_d59_47;
	wire [WIDTH-1:0] wire_d59_48;
	wire [WIDTH-1:0] wire_d59_49;
	wire [WIDTH-1:0] wire_d59_50;
	wire [WIDTH-1:0] wire_d59_51;
	wire [WIDTH-1:0] wire_d59_52;
	wire [WIDTH-1:0] wire_d59_53;
	wire [WIDTH-1:0] wire_d59_54;
	wire [WIDTH-1:0] wire_d59_55;
	wire [WIDTH-1:0] wire_d59_56;
	wire [WIDTH-1:0] wire_d59_57;
	wire [WIDTH-1:0] wire_d59_58;
	wire [WIDTH-1:0] wire_d59_59;
	wire [WIDTH-1:0] wire_d59_60;
	wire [WIDTH-1:0] wire_d59_61;
	wire [WIDTH-1:0] wire_d59_62;
	wire [WIDTH-1:0] wire_d59_63;
	wire [WIDTH-1:0] wire_d59_64;
	wire [WIDTH-1:0] wire_d59_65;
	wire [WIDTH-1:0] wire_d59_66;
	wire [WIDTH-1:0] wire_d59_67;
	wire [WIDTH-1:0] wire_d59_68;
	wire [WIDTH-1:0] wire_d59_69;
	wire [WIDTH-1:0] wire_d59_70;
	wire [WIDTH-1:0] wire_d59_71;
	wire [WIDTH-1:0] wire_d59_72;
	wire [WIDTH-1:0] wire_d59_73;
	wire [WIDTH-1:0] wire_d59_74;
	wire [WIDTH-1:0] wire_d59_75;
	wire [WIDTH-1:0] wire_d59_76;
	wire [WIDTH-1:0] wire_d59_77;
	wire [WIDTH-1:0] wire_d59_78;

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance101(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance102(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance103(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance104(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance105(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance106(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance107(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance108(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance109(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1029(.data_in(wire_d0_28),.data_out(wire_d0_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1030(.data_in(wire_d0_29),.data_out(wire_d0_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1031(.data_in(wire_d0_30),.data_out(wire_d0_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1032(.data_in(wire_d0_31),.data_out(wire_d0_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1033(.data_in(wire_d0_32),.data_out(wire_d0_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1034(.data_in(wire_d0_33),.data_out(wire_d0_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1035(.data_in(wire_d0_34),.data_out(wire_d0_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1036(.data_in(wire_d0_35),.data_out(wire_d0_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1037(.data_in(wire_d0_36),.data_out(wire_d0_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1038(.data_in(wire_d0_37),.data_out(wire_d0_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1039(.data_in(wire_d0_38),.data_out(wire_d0_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1040(.data_in(wire_d0_39),.data_out(wire_d0_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1041(.data_in(wire_d0_40),.data_out(wire_d0_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1042(.data_in(wire_d0_41),.data_out(wire_d0_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1043(.data_in(wire_d0_42),.data_out(wire_d0_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1044(.data_in(wire_d0_43),.data_out(wire_d0_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1045(.data_in(wire_d0_44),.data_out(wire_d0_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1046(.data_in(wire_d0_45),.data_out(wire_d0_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1047(.data_in(wire_d0_46),.data_out(wire_d0_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1048(.data_in(wire_d0_47),.data_out(wire_d0_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1049(.data_in(wire_d0_48),.data_out(wire_d0_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1050(.data_in(wire_d0_49),.data_out(wire_d0_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1051(.data_in(wire_d0_50),.data_out(wire_d0_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1052(.data_in(wire_d0_51),.data_out(wire_d0_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1053(.data_in(wire_d0_52),.data_out(wire_d0_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1054(.data_in(wire_d0_53),.data_out(wire_d0_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1055(.data_in(wire_d0_54),.data_out(wire_d0_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1056(.data_in(wire_d0_55),.data_out(wire_d0_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1057(.data_in(wire_d0_56),.data_out(wire_d0_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1058(.data_in(wire_d0_57),.data_out(wire_d0_58),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1059(.data_in(wire_d0_58),.data_out(wire_d0_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1060(.data_in(wire_d0_59),.data_out(wire_d0_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1061(.data_in(wire_d0_60),.data_out(wire_d0_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1062(.data_in(wire_d0_61),.data_out(wire_d0_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1063(.data_in(wire_d0_62),.data_out(wire_d0_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1064(.data_in(wire_d0_63),.data_out(wire_d0_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1065(.data_in(wire_d0_64),.data_out(wire_d0_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1066(.data_in(wire_d0_65),.data_out(wire_d0_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1067(.data_in(wire_d0_66),.data_out(wire_d0_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1068(.data_in(wire_d0_67),.data_out(wire_d0_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1069(.data_in(wire_d0_68),.data_out(wire_d0_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1070(.data_in(wire_d0_69),.data_out(wire_d0_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1071(.data_in(wire_d0_70),.data_out(wire_d0_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1072(.data_in(wire_d0_71),.data_out(wire_d0_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1073(.data_in(wire_d0_72),.data_out(wire_d0_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1074(.data_in(wire_d0_73),.data_out(wire_d0_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1075(.data_in(wire_d0_74),.data_out(wire_d0_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1076(.data_in(wire_d0_75),.data_out(wire_d0_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1077(.data_in(wire_d0_76),.data_out(wire_d0_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1078(.data_in(wire_d0_77),.data_out(wire_d0_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1079(.data_in(wire_d0_78),.data_out(d_out0),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance210(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance211(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance213(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance214(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance215(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance216(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance217(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance218(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance219(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2129(.data_in(wire_d1_28),.data_out(wire_d1_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2130(.data_in(wire_d1_29),.data_out(wire_d1_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2131(.data_in(wire_d1_30),.data_out(wire_d1_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2132(.data_in(wire_d1_31),.data_out(wire_d1_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2133(.data_in(wire_d1_32),.data_out(wire_d1_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2134(.data_in(wire_d1_33),.data_out(wire_d1_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2135(.data_in(wire_d1_34),.data_out(wire_d1_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2136(.data_in(wire_d1_35),.data_out(wire_d1_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2137(.data_in(wire_d1_36),.data_out(wire_d1_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2138(.data_in(wire_d1_37),.data_out(wire_d1_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2139(.data_in(wire_d1_38),.data_out(wire_d1_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2140(.data_in(wire_d1_39),.data_out(wire_d1_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2141(.data_in(wire_d1_40),.data_out(wire_d1_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2142(.data_in(wire_d1_41),.data_out(wire_d1_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2143(.data_in(wire_d1_42),.data_out(wire_d1_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2144(.data_in(wire_d1_43),.data_out(wire_d1_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2145(.data_in(wire_d1_44),.data_out(wire_d1_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2146(.data_in(wire_d1_45),.data_out(wire_d1_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2147(.data_in(wire_d1_46),.data_out(wire_d1_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2148(.data_in(wire_d1_47),.data_out(wire_d1_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2149(.data_in(wire_d1_48),.data_out(wire_d1_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2150(.data_in(wire_d1_49),.data_out(wire_d1_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2151(.data_in(wire_d1_50),.data_out(wire_d1_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2152(.data_in(wire_d1_51),.data_out(wire_d1_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2153(.data_in(wire_d1_52),.data_out(wire_d1_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2154(.data_in(wire_d1_53),.data_out(wire_d1_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2155(.data_in(wire_d1_54),.data_out(wire_d1_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2156(.data_in(wire_d1_55),.data_out(wire_d1_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2157(.data_in(wire_d1_56),.data_out(wire_d1_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2158(.data_in(wire_d1_57),.data_out(wire_d1_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2159(.data_in(wire_d1_58),.data_out(wire_d1_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2160(.data_in(wire_d1_59),.data_out(wire_d1_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2161(.data_in(wire_d1_60),.data_out(wire_d1_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2162(.data_in(wire_d1_61),.data_out(wire_d1_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2163(.data_in(wire_d1_62),.data_out(wire_d1_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2164(.data_in(wire_d1_63),.data_out(wire_d1_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2165(.data_in(wire_d1_64),.data_out(wire_d1_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2166(.data_in(wire_d1_65),.data_out(wire_d1_66),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2167(.data_in(wire_d1_66),.data_out(wire_d1_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2168(.data_in(wire_d1_67),.data_out(wire_d1_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2169(.data_in(wire_d1_68),.data_out(wire_d1_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2170(.data_in(wire_d1_69),.data_out(wire_d1_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2171(.data_in(wire_d1_70),.data_out(wire_d1_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2172(.data_in(wire_d1_71),.data_out(wire_d1_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2173(.data_in(wire_d1_72),.data_out(wire_d1_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2174(.data_in(wire_d1_73),.data_out(wire_d1_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2175(.data_in(wire_d1_74),.data_out(wire_d1_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2176(.data_in(wire_d1_75),.data_out(wire_d1_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2177(.data_in(wire_d1_76),.data_out(wire_d1_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2178(.data_in(wire_d1_77),.data_out(wire_d1_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2179(.data_in(wire_d1_78),.data_out(d_out1),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance320(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance321(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance322(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance324(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance325(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance326(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance327(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance328(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance329(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3229(.data_in(wire_d2_28),.data_out(wire_d2_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3230(.data_in(wire_d2_29),.data_out(wire_d2_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3231(.data_in(wire_d2_30),.data_out(wire_d2_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3232(.data_in(wire_d2_31),.data_out(wire_d2_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3233(.data_in(wire_d2_32),.data_out(wire_d2_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3234(.data_in(wire_d2_33),.data_out(wire_d2_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3235(.data_in(wire_d2_34),.data_out(wire_d2_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3236(.data_in(wire_d2_35),.data_out(wire_d2_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3237(.data_in(wire_d2_36),.data_out(wire_d2_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3238(.data_in(wire_d2_37),.data_out(wire_d2_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3239(.data_in(wire_d2_38),.data_out(wire_d2_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3240(.data_in(wire_d2_39),.data_out(wire_d2_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3241(.data_in(wire_d2_40),.data_out(wire_d2_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3242(.data_in(wire_d2_41),.data_out(wire_d2_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3243(.data_in(wire_d2_42),.data_out(wire_d2_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3244(.data_in(wire_d2_43),.data_out(wire_d2_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3245(.data_in(wire_d2_44),.data_out(wire_d2_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3246(.data_in(wire_d2_45),.data_out(wire_d2_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3247(.data_in(wire_d2_46),.data_out(wire_d2_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3248(.data_in(wire_d2_47),.data_out(wire_d2_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3249(.data_in(wire_d2_48),.data_out(wire_d2_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3250(.data_in(wire_d2_49),.data_out(wire_d2_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3251(.data_in(wire_d2_50),.data_out(wire_d2_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3252(.data_in(wire_d2_51),.data_out(wire_d2_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3253(.data_in(wire_d2_52),.data_out(wire_d2_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3254(.data_in(wire_d2_53),.data_out(wire_d2_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3255(.data_in(wire_d2_54),.data_out(wire_d2_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3256(.data_in(wire_d2_55),.data_out(wire_d2_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3257(.data_in(wire_d2_56),.data_out(wire_d2_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3258(.data_in(wire_d2_57),.data_out(wire_d2_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3259(.data_in(wire_d2_58),.data_out(wire_d2_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3260(.data_in(wire_d2_59),.data_out(wire_d2_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3261(.data_in(wire_d2_60),.data_out(wire_d2_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3262(.data_in(wire_d2_61),.data_out(wire_d2_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3263(.data_in(wire_d2_62),.data_out(wire_d2_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3264(.data_in(wire_d2_63),.data_out(wire_d2_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3265(.data_in(wire_d2_64),.data_out(wire_d2_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3266(.data_in(wire_d2_65),.data_out(wire_d2_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3267(.data_in(wire_d2_66),.data_out(wire_d2_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3268(.data_in(wire_d2_67),.data_out(wire_d2_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3269(.data_in(wire_d2_68),.data_out(wire_d2_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3270(.data_in(wire_d2_69),.data_out(wire_d2_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3271(.data_in(wire_d2_70),.data_out(wire_d2_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3272(.data_in(wire_d2_71),.data_out(wire_d2_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3273(.data_in(wire_d2_72),.data_out(wire_d2_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3274(.data_in(wire_d2_73),.data_out(wire_d2_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3275(.data_in(wire_d2_74),.data_out(wire_d2_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3276(.data_in(wire_d2_75),.data_out(wire_d2_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3277(.data_in(wire_d2_76),.data_out(wire_d2_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3278(.data_in(wire_d2_77),.data_out(wire_d2_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3279(.data_in(wire_d2_78),.data_out(d_out2),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance430(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance431(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance432(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance433(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance434(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance435(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance436(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance437(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance438(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance439(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4329(.data_in(wire_d3_28),.data_out(wire_d3_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4330(.data_in(wire_d3_29),.data_out(wire_d3_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4331(.data_in(wire_d3_30),.data_out(wire_d3_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4332(.data_in(wire_d3_31),.data_out(wire_d3_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4333(.data_in(wire_d3_32),.data_out(wire_d3_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4334(.data_in(wire_d3_33),.data_out(wire_d3_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4335(.data_in(wire_d3_34),.data_out(wire_d3_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4336(.data_in(wire_d3_35),.data_out(wire_d3_36),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4337(.data_in(wire_d3_36),.data_out(wire_d3_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4338(.data_in(wire_d3_37),.data_out(wire_d3_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4339(.data_in(wire_d3_38),.data_out(wire_d3_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4340(.data_in(wire_d3_39),.data_out(wire_d3_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4341(.data_in(wire_d3_40),.data_out(wire_d3_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4342(.data_in(wire_d3_41),.data_out(wire_d3_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4343(.data_in(wire_d3_42),.data_out(wire_d3_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4344(.data_in(wire_d3_43),.data_out(wire_d3_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4345(.data_in(wire_d3_44),.data_out(wire_d3_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4346(.data_in(wire_d3_45),.data_out(wire_d3_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4347(.data_in(wire_d3_46),.data_out(wire_d3_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4348(.data_in(wire_d3_47),.data_out(wire_d3_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4349(.data_in(wire_d3_48),.data_out(wire_d3_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4350(.data_in(wire_d3_49),.data_out(wire_d3_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4351(.data_in(wire_d3_50),.data_out(wire_d3_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4352(.data_in(wire_d3_51),.data_out(wire_d3_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4353(.data_in(wire_d3_52),.data_out(wire_d3_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4354(.data_in(wire_d3_53),.data_out(wire_d3_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4355(.data_in(wire_d3_54),.data_out(wire_d3_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4356(.data_in(wire_d3_55),.data_out(wire_d3_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4357(.data_in(wire_d3_56),.data_out(wire_d3_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4358(.data_in(wire_d3_57),.data_out(wire_d3_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4359(.data_in(wire_d3_58),.data_out(wire_d3_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4360(.data_in(wire_d3_59),.data_out(wire_d3_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4361(.data_in(wire_d3_60),.data_out(wire_d3_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4362(.data_in(wire_d3_61),.data_out(wire_d3_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4363(.data_in(wire_d3_62),.data_out(wire_d3_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4364(.data_in(wire_d3_63),.data_out(wire_d3_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4365(.data_in(wire_d3_64),.data_out(wire_d3_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4366(.data_in(wire_d3_65),.data_out(wire_d3_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4367(.data_in(wire_d3_66),.data_out(wire_d3_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4368(.data_in(wire_d3_67),.data_out(wire_d3_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4369(.data_in(wire_d3_68),.data_out(wire_d3_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4370(.data_in(wire_d3_69),.data_out(wire_d3_70),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4371(.data_in(wire_d3_70),.data_out(wire_d3_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4372(.data_in(wire_d3_71),.data_out(wire_d3_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4373(.data_in(wire_d3_72),.data_out(wire_d3_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4374(.data_in(wire_d3_73),.data_out(wire_d3_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4375(.data_in(wire_d3_74),.data_out(wire_d3_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4376(.data_in(wire_d3_75),.data_out(wire_d3_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4377(.data_in(wire_d3_76),.data_out(wire_d3_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4378(.data_in(wire_d3_77),.data_out(wire_d3_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4379(.data_in(wire_d3_78),.data_out(d_out3),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance540(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance541(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance542(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance543(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance544(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance545(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance546(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance547(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance548(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance549(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5429(.data_in(wire_d4_28),.data_out(wire_d4_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5430(.data_in(wire_d4_29),.data_out(wire_d4_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5431(.data_in(wire_d4_30),.data_out(wire_d4_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5432(.data_in(wire_d4_31),.data_out(wire_d4_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5433(.data_in(wire_d4_32),.data_out(wire_d4_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5434(.data_in(wire_d4_33),.data_out(wire_d4_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5435(.data_in(wire_d4_34),.data_out(wire_d4_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5436(.data_in(wire_d4_35),.data_out(wire_d4_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5437(.data_in(wire_d4_36),.data_out(wire_d4_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5438(.data_in(wire_d4_37),.data_out(wire_d4_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5439(.data_in(wire_d4_38),.data_out(wire_d4_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5440(.data_in(wire_d4_39),.data_out(wire_d4_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5441(.data_in(wire_d4_40),.data_out(wire_d4_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5442(.data_in(wire_d4_41),.data_out(wire_d4_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5443(.data_in(wire_d4_42),.data_out(wire_d4_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5444(.data_in(wire_d4_43),.data_out(wire_d4_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5445(.data_in(wire_d4_44),.data_out(wire_d4_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5446(.data_in(wire_d4_45),.data_out(wire_d4_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5447(.data_in(wire_d4_46),.data_out(wire_d4_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5448(.data_in(wire_d4_47),.data_out(wire_d4_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5449(.data_in(wire_d4_48),.data_out(wire_d4_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5450(.data_in(wire_d4_49),.data_out(wire_d4_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5451(.data_in(wire_d4_50),.data_out(wire_d4_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5452(.data_in(wire_d4_51),.data_out(wire_d4_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5453(.data_in(wire_d4_52),.data_out(wire_d4_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5454(.data_in(wire_d4_53),.data_out(wire_d4_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5455(.data_in(wire_d4_54),.data_out(wire_d4_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5456(.data_in(wire_d4_55),.data_out(wire_d4_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5457(.data_in(wire_d4_56),.data_out(wire_d4_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5458(.data_in(wire_d4_57),.data_out(wire_d4_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5459(.data_in(wire_d4_58),.data_out(wire_d4_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5460(.data_in(wire_d4_59),.data_out(wire_d4_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5461(.data_in(wire_d4_60),.data_out(wire_d4_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5462(.data_in(wire_d4_61),.data_out(wire_d4_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5463(.data_in(wire_d4_62),.data_out(wire_d4_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5464(.data_in(wire_d4_63),.data_out(wire_d4_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5465(.data_in(wire_d4_64),.data_out(wire_d4_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5466(.data_in(wire_d4_65),.data_out(wire_d4_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5467(.data_in(wire_d4_66),.data_out(wire_d4_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5468(.data_in(wire_d4_67),.data_out(wire_d4_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5469(.data_in(wire_d4_68),.data_out(wire_d4_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5470(.data_in(wire_d4_69),.data_out(wire_d4_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5471(.data_in(wire_d4_70),.data_out(wire_d4_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5472(.data_in(wire_d4_71),.data_out(wire_d4_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5473(.data_in(wire_d4_72),.data_out(wire_d4_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5474(.data_in(wire_d4_73),.data_out(wire_d4_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5475(.data_in(wire_d4_74),.data_out(wire_d4_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5476(.data_in(wire_d4_75),.data_out(wire_d4_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5477(.data_in(wire_d4_76),.data_out(wire_d4_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5478(.data_in(wire_d4_77),.data_out(wire_d4_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5479(.data_in(wire_d4_78),.data_out(d_out4),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance650(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	invertion #(.WIDTH(WIDTH)) invertion_instance651(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance652(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance653(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance654(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance655(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance656(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance657(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance658(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance659(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6529(.data_in(wire_d5_28),.data_out(wire_d5_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6530(.data_in(wire_d5_29),.data_out(wire_d5_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6531(.data_in(wire_d5_30),.data_out(wire_d5_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6532(.data_in(wire_d5_31),.data_out(wire_d5_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6533(.data_in(wire_d5_32),.data_out(wire_d5_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6534(.data_in(wire_d5_33),.data_out(wire_d5_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6535(.data_in(wire_d5_34),.data_out(wire_d5_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6536(.data_in(wire_d5_35),.data_out(wire_d5_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6537(.data_in(wire_d5_36),.data_out(wire_d5_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6538(.data_in(wire_d5_37),.data_out(wire_d5_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6539(.data_in(wire_d5_38),.data_out(wire_d5_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6540(.data_in(wire_d5_39),.data_out(wire_d5_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6541(.data_in(wire_d5_40),.data_out(wire_d5_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6542(.data_in(wire_d5_41),.data_out(wire_d5_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6543(.data_in(wire_d5_42),.data_out(wire_d5_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6544(.data_in(wire_d5_43),.data_out(wire_d5_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6545(.data_in(wire_d5_44),.data_out(wire_d5_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6546(.data_in(wire_d5_45),.data_out(wire_d5_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6547(.data_in(wire_d5_46),.data_out(wire_d5_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6548(.data_in(wire_d5_47),.data_out(wire_d5_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6549(.data_in(wire_d5_48),.data_out(wire_d5_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6550(.data_in(wire_d5_49),.data_out(wire_d5_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6551(.data_in(wire_d5_50),.data_out(wire_d5_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6552(.data_in(wire_d5_51),.data_out(wire_d5_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6553(.data_in(wire_d5_52),.data_out(wire_d5_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6554(.data_in(wire_d5_53),.data_out(wire_d5_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6555(.data_in(wire_d5_54),.data_out(wire_d5_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6556(.data_in(wire_d5_55),.data_out(wire_d5_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6557(.data_in(wire_d5_56),.data_out(wire_d5_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6558(.data_in(wire_d5_57),.data_out(wire_d5_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6559(.data_in(wire_d5_58),.data_out(wire_d5_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6560(.data_in(wire_d5_59),.data_out(wire_d5_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6561(.data_in(wire_d5_60),.data_out(wire_d5_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6562(.data_in(wire_d5_61),.data_out(wire_d5_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6563(.data_in(wire_d5_62),.data_out(wire_d5_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6564(.data_in(wire_d5_63),.data_out(wire_d5_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6565(.data_in(wire_d5_64),.data_out(wire_d5_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6566(.data_in(wire_d5_65),.data_out(wire_d5_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6567(.data_in(wire_d5_66),.data_out(wire_d5_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6568(.data_in(wire_d5_67),.data_out(wire_d5_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6569(.data_in(wire_d5_68),.data_out(wire_d5_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6570(.data_in(wire_d5_69),.data_out(wire_d5_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6571(.data_in(wire_d5_70),.data_out(wire_d5_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6572(.data_in(wire_d5_71),.data_out(wire_d5_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6573(.data_in(wire_d5_72),.data_out(wire_d5_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6574(.data_in(wire_d5_73),.data_out(wire_d5_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6575(.data_in(wire_d5_74),.data_out(wire_d5_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6576(.data_in(wire_d5_75),.data_out(wire_d5_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6577(.data_in(wire_d5_76),.data_out(wire_d5_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6578(.data_in(wire_d5_77),.data_out(wire_d5_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6579(.data_in(wire_d5_78),.data_out(d_out5),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance760(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	large_mux #(.WIDTH(WIDTH)) large_mux_instance761(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance762(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance763(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance764(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance765(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance766(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance768(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance769(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7629(.data_in(wire_d6_28),.data_out(wire_d6_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7630(.data_in(wire_d6_29),.data_out(wire_d6_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7631(.data_in(wire_d6_30),.data_out(wire_d6_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7632(.data_in(wire_d6_31),.data_out(wire_d6_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7633(.data_in(wire_d6_32),.data_out(wire_d6_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7634(.data_in(wire_d6_33),.data_out(wire_d6_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7635(.data_in(wire_d6_34),.data_out(wire_d6_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7636(.data_in(wire_d6_35),.data_out(wire_d6_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7637(.data_in(wire_d6_36),.data_out(wire_d6_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7638(.data_in(wire_d6_37),.data_out(wire_d6_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7639(.data_in(wire_d6_38),.data_out(wire_d6_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7640(.data_in(wire_d6_39),.data_out(wire_d6_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7641(.data_in(wire_d6_40),.data_out(wire_d6_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7642(.data_in(wire_d6_41),.data_out(wire_d6_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7643(.data_in(wire_d6_42),.data_out(wire_d6_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7644(.data_in(wire_d6_43),.data_out(wire_d6_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7645(.data_in(wire_d6_44),.data_out(wire_d6_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7646(.data_in(wire_d6_45),.data_out(wire_d6_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7647(.data_in(wire_d6_46),.data_out(wire_d6_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7648(.data_in(wire_d6_47),.data_out(wire_d6_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7649(.data_in(wire_d6_48),.data_out(wire_d6_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7650(.data_in(wire_d6_49),.data_out(wire_d6_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7651(.data_in(wire_d6_50),.data_out(wire_d6_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7652(.data_in(wire_d6_51),.data_out(wire_d6_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7653(.data_in(wire_d6_52),.data_out(wire_d6_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7654(.data_in(wire_d6_53),.data_out(wire_d6_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7655(.data_in(wire_d6_54),.data_out(wire_d6_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7656(.data_in(wire_d6_55),.data_out(wire_d6_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7657(.data_in(wire_d6_56),.data_out(wire_d6_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7658(.data_in(wire_d6_57),.data_out(wire_d6_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7659(.data_in(wire_d6_58),.data_out(wire_d6_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7660(.data_in(wire_d6_59),.data_out(wire_d6_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7661(.data_in(wire_d6_60),.data_out(wire_d6_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7662(.data_in(wire_d6_61),.data_out(wire_d6_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7663(.data_in(wire_d6_62),.data_out(wire_d6_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7664(.data_in(wire_d6_63),.data_out(wire_d6_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7665(.data_in(wire_d6_64),.data_out(wire_d6_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7666(.data_in(wire_d6_65),.data_out(wire_d6_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7667(.data_in(wire_d6_66),.data_out(wire_d6_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7668(.data_in(wire_d6_67),.data_out(wire_d6_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7669(.data_in(wire_d6_68),.data_out(wire_d6_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7670(.data_in(wire_d6_69),.data_out(wire_d6_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7671(.data_in(wire_d6_70),.data_out(wire_d6_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7672(.data_in(wire_d6_71),.data_out(wire_d6_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7673(.data_in(wire_d6_72),.data_out(wire_d6_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7674(.data_in(wire_d6_73),.data_out(wire_d6_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7675(.data_in(wire_d6_74),.data_out(wire_d6_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7676(.data_in(wire_d6_75),.data_out(wire_d6_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7677(.data_in(wire_d6_76),.data_out(wire_d6_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7678(.data_in(wire_d6_77),.data_out(wire_d6_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7679(.data_in(wire_d6_78),.data_out(d_out6),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance870(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance871(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance872(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance873(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance874(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance875(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance876(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance877(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance878(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance879(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8729(.data_in(wire_d7_28),.data_out(wire_d7_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8730(.data_in(wire_d7_29),.data_out(wire_d7_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8731(.data_in(wire_d7_30),.data_out(wire_d7_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8732(.data_in(wire_d7_31),.data_out(wire_d7_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8733(.data_in(wire_d7_32),.data_out(wire_d7_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8734(.data_in(wire_d7_33),.data_out(wire_d7_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8735(.data_in(wire_d7_34),.data_out(wire_d7_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8736(.data_in(wire_d7_35),.data_out(wire_d7_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8737(.data_in(wire_d7_36),.data_out(wire_d7_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8738(.data_in(wire_d7_37),.data_out(wire_d7_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8739(.data_in(wire_d7_38),.data_out(wire_d7_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8740(.data_in(wire_d7_39),.data_out(wire_d7_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8741(.data_in(wire_d7_40),.data_out(wire_d7_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8742(.data_in(wire_d7_41),.data_out(wire_d7_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8743(.data_in(wire_d7_42),.data_out(wire_d7_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8744(.data_in(wire_d7_43),.data_out(wire_d7_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8745(.data_in(wire_d7_44),.data_out(wire_d7_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8746(.data_in(wire_d7_45),.data_out(wire_d7_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8747(.data_in(wire_d7_46),.data_out(wire_d7_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8748(.data_in(wire_d7_47),.data_out(wire_d7_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8749(.data_in(wire_d7_48),.data_out(wire_d7_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8750(.data_in(wire_d7_49),.data_out(wire_d7_50),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8751(.data_in(wire_d7_50),.data_out(wire_d7_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8752(.data_in(wire_d7_51),.data_out(wire_d7_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8753(.data_in(wire_d7_52),.data_out(wire_d7_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8754(.data_in(wire_d7_53),.data_out(wire_d7_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8755(.data_in(wire_d7_54),.data_out(wire_d7_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8756(.data_in(wire_d7_55),.data_out(wire_d7_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8757(.data_in(wire_d7_56),.data_out(wire_d7_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8758(.data_in(wire_d7_57),.data_out(wire_d7_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8759(.data_in(wire_d7_58),.data_out(wire_d7_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8760(.data_in(wire_d7_59),.data_out(wire_d7_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8761(.data_in(wire_d7_60),.data_out(wire_d7_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8762(.data_in(wire_d7_61),.data_out(wire_d7_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8763(.data_in(wire_d7_62),.data_out(wire_d7_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8764(.data_in(wire_d7_63),.data_out(wire_d7_64),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8765(.data_in(wire_d7_64),.data_out(wire_d7_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8766(.data_in(wire_d7_65),.data_out(wire_d7_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8767(.data_in(wire_d7_66),.data_out(wire_d7_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8768(.data_in(wire_d7_67),.data_out(wire_d7_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8769(.data_in(wire_d7_68),.data_out(wire_d7_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8770(.data_in(wire_d7_69),.data_out(wire_d7_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8771(.data_in(wire_d7_70),.data_out(wire_d7_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8772(.data_in(wire_d7_71),.data_out(wire_d7_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8773(.data_in(wire_d7_72),.data_out(wire_d7_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8774(.data_in(wire_d7_73),.data_out(wire_d7_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8775(.data_in(wire_d7_74),.data_out(wire_d7_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8776(.data_in(wire_d7_75),.data_out(wire_d7_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8777(.data_in(wire_d7_76),.data_out(wire_d7_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8778(.data_in(wire_d7_77),.data_out(wire_d7_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8779(.data_in(wire_d7_78),.data_out(d_out7),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance980(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	decoder_top #(.WIDTH(WIDTH)) decoder_instance981(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance982(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance983(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance984(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance985(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance986(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance987(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance988(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance989(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9829(.data_in(wire_d8_28),.data_out(wire_d8_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9830(.data_in(wire_d8_29),.data_out(wire_d8_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9831(.data_in(wire_d8_30),.data_out(wire_d8_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9832(.data_in(wire_d8_31),.data_out(wire_d8_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9833(.data_in(wire_d8_32),.data_out(wire_d8_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9834(.data_in(wire_d8_33),.data_out(wire_d8_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9835(.data_in(wire_d8_34),.data_out(wire_d8_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9836(.data_in(wire_d8_35),.data_out(wire_d8_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9837(.data_in(wire_d8_36),.data_out(wire_d8_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9838(.data_in(wire_d8_37),.data_out(wire_d8_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9839(.data_in(wire_d8_38),.data_out(wire_d8_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9840(.data_in(wire_d8_39),.data_out(wire_d8_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9841(.data_in(wire_d8_40),.data_out(wire_d8_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9842(.data_in(wire_d8_41),.data_out(wire_d8_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9843(.data_in(wire_d8_42),.data_out(wire_d8_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9844(.data_in(wire_d8_43),.data_out(wire_d8_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9845(.data_in(wire_d8_44),.data_out(wire_d8_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9846(.data_in(wire_d8_45),.data_out(wire_d8_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9847(.data_in(wire_d8_46),.data_out(wire_d8_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9848(.data_in(wire_d8_47),.data_out(wire_d8_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9849(.data_in(wire_d8_48),.data_out(wire_d8_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9850(.data_in(wire_d8_49),.data_out(wire_d8_50),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9851(.data_in(wire_d8_50),.data_out(wire_d8_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9852(.data_in(wire_d8_51),.data_out(wire_d8_52),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9853(.data_in(wire_d8_52),.data_out(wire_d8_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9854(.data_in(wire_d8_53),.data_out(wire_d8_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9855(.data_in(wire_d8_54),.data_out(wire_d8_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9856(.data_in(wire_d8_55),.data_out(wire_d8_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9857(.data_in(wire_d8_56),.data_out(wire_d8_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9858(.data_in(wire_d8_57),.data_out(wire_d8_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9859(.data_in(wire_d8_58),.data_out(wire_d8_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9860(.data_in(wire_d8_59),.data_out(wire_d8_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9861(.data_in(wire_d8_60),.data_out(wire_d8_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9862(.data_in(wire_d8_61),.data_out(wire_d8_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9863(.data_in(wire_d8_62),.data_out(wire_d8_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9864(.data_in(wire_d8_63),.data_out(wire_d8_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9865(.data_in(wire_d8_64),.data_out(wire_d8_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9866(.data_in(wire_d8_65),.data_out(wire_d8_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9867(.data_in(wire_d8_66),.data_out(wire_d8_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9868(.data_in(wire_d8_67),.data_out(wire_d8_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9869(.data_in(wire_d8_68),.data_out(wire_d8_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9870(.data_in(wire_d8_69),.data_out(wire_d8_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9871(.data_in(wire_d8_70),.data_out(wire_d8_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9872(.data_in(wire_d8_71),.data_out(wire_d8_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9873(.data_in(wire_d8_72),.data_out(wire_d8_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9874(.data_in(wire_d8_73),.data_out(wire_d8_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9875(.data_in(wire_d8_74),.data_out(wire_d8_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9876(.data_in(wire_d8_75),.data_out(wire_d8_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9877(.data_in(wire_d8_76),.data_out(wire_d8_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9878(.data_in(wire_d8_77),.data_out(wire_d8_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9879(.data_in(wire_d8_78),.data_out(d_out8),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance10090(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10091(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10092(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10093(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10094(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10095(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10096(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10097(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10098(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10099(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100929(.data_in(wire_d9_28),.data_out(wire_d9_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100930(.data_in(wire_d9_29),.data_out(wire_d9_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100931(.data_in(wire_d9_30),.data_out(wire_d9_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100932(.data_in(wire_d9_31),.data_out(wire_d9_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100933(.data_in(wire_d9_32),.data_out(wire_d9_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100934(.data_in(wire_d9_33),.data_out(wire_d9_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100935(.data_in(wire_d9_34),.data_out(wire_d9_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100936(.data_in(wire_d9_35),.data_out(wire_d9_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100937(.data_in(wire_d9_36),.data_out(wire_d9_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100938(.data_in(wire_d9_37),.data_out(wire_d9_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100939(.data_in(wire_d9_38),.data_out(wire_d9_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100940(.data_in(wire_d9_39),.data_out(wire_d9_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100941(.data_in(wire_d9_40),.data_out(wire_d9_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100942(.data_in(wire_d9_41),.data_out(wire_d9_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100943(.data_in(wire_d9_42),.data_out(wire_d9_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100944(.data_in(wire_d9_43),.data_out(wire_d9_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100945(.data_in(wire_d9_44),.data_out(wire_d9_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100946(.data_in(wire_d9_45),.data_out(wire_d9_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100947(.data_in(wire_d9_46),.data_out(wire_d9_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100948(.data_in(wire_d9_47),.data_out(wire_d9_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100949(.data_in(wire_d9_48),.data_out(wire_d9_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100950(.data_in(wire_d9_49),.data_out(wire_d9_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100951(.data_in(wire_d9_50),.data_out(wire_d9_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100952(.data_in(wire_d9_51),.data_out(wire_d9_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100953(.data_in(wire_d9_52),.data_out(wire_d9_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100954(.data_in(wire_d9_53),.data_out(wire_d9_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100955(.data_in(wire_d9_54),.data_out(wire_d9_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100956(.data_in(wire_d9_55),.data_out(wire_d9_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100957(.data_in(wire_d9_56),.data_out(wire_d9_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100958(.data_in(wire_d9_57),.data_out(wire_d9_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100959(.data_in(wire_d9_58),.data_out(wire_d9_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100960(.data_in(wire_d9_59),.data_out(wire_d9_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100961(.data_in(wire_d9_60),.data_out(wire_d9_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100962(.data_in(wire_d9_61),.data_out(wire_d9_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100963(.data_in(wire_d9_62),.data_out(wire_d9_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100964(.data_in(wire_d9_63),.data_out(wire_d9_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100965(.data_in(wire_d9_64),.data_out(wire_d9_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100966(.data_in(wire_d9_65),.data_out(wire_d9_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100967(.data_in(wire_d9_66),.data_out(wire_d9_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100968(.data_in(wire_d9_67),.data_out(wire_d9_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100969(.data_in(wire_d9_68),.data_out(wire_d9_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100970(.data_in(wire_d9_69),.data_out(wire_d9_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100971(.data_in(wire_d9_70),.data_out(wire_d9_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100972(.data_in(wire_d9_71),.data_out(wire_d9_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100973(.data_in(wire_d9_72),.data_out(wire_d9_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100974(.data_in(wire_d9_73),.data_out(wire_d9_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100975(.data_in(wire_d9_74),.data_out(wire_d9_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100976(.data_in(wire_d9_75),.data_out(wire_d9_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100977(.data_in(wire_d9_76),.data_out(wire_d9_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100978(.data_in(wire_d9_77),.data_out(wire_d9_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100979(.data_in(wire_d9_78),.data_out(d_out9),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance110100(.data_in(d_in10),.data_out(wire_d10_0),.clk(clk),.rst(rst));            //channel 11
	large_mux #(.WIDTH(WIDTH)) large_mux_instance110101(.data_in(wire_d10_0),.data_out(wire_d10_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance110102(.data_in(wire_d10_1),.data_out(wire_d10_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance110103(.data_in(wire_d10_2),.data_out(wire_d10_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance110104(.data_in(wire_d10_3),.data_out(wire_d10_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance110105(.data_in(wire_d10_4),.data_out(wire_d10_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance110106(.data_in(wire_d10_5),.data_out(wire_d10_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance110107(.data_in(wire_d10_6),.data_out(wire_d10_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance110108(.data_in(wire_d10_7),.data_out(wire_d10_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance110109(.data_in(wire_d10_8),.data_out(wire_d10_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101010(.data_in(wire_d10_9),.data_out(wire_d10_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101011(.data_in(wire_d10_10),.data_out(wire_d10_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101012(.data_in(wire_d10_11),.data_out(wire_d10_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101013(.data_in(wire_d10_12),.data_out(wire_d10_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101014(.data_in(wire_d10_13),.data_out(wire_d10_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101015(.data_in(wire_d10_14),.data_out(wire_d10_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101016(.data_in(wire_d10_15),.data_out(wire_d10_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101017(.data_in(wire_d10_16),.data_out(wire_d10_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101018(.data_in(wire_d10_17),.data_out(wire_d10_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101019(.data_in(wire_d10_18),.data_out(wire_d10_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101020(.data_in(wire_d10_19),.data_out(wire_d10_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101021(.data_in(wire_d10_20),.data_out(wire_d10_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101022(.data_in(wire_d10_21),.data_out(wire_d10_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101023(.data_in(wire_d10_22),.data_out(wire_d10_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101024(.data_in(wire_d10_23),.data_out(wire_d10_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101025(.data_in(wire_d10_24),.data_out(wire_d10_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101026(.data_in(wire_d10_25),.data_out(wire_d10_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101027(.data_in(wire_d10_26),.data_out(wire_d10_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101028(.data_in(wire_d10_27),.data_out(wire_d10_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101029(.data_in(wire_d10_28),.data_out(wire_d10_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101030(.data_in(wire_d10_29),.data_out(wire_d10_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101031(.data_in(wire_d10_30),.data_out(wire_d10_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101032(.data_in(wire_d10_31),.data_out(wire_d10_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101033(.data_in(wire_d10_32),.data_out(wire_d10_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101034(.data_in(wire_d10_33),.data_out(wire_d10_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101035(.data_in(wire_d10_34),.data_out(wire_d10_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101036(.data_in(wire_d10_35),.data_out(wire_d10_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101037(.data_in(wire_d10_36),.data_out(wire_d10_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101038(.data_in(wire_d10_37),.data_out(wire_d10_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101039(.data_in(wire_d10_38),.data_out(wire_d10_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101040(.data_in(wire_d10_39),.data_out(wire_d10_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101041(.data_in(wire_d10_40),.data_out(wire_d10_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101042(.data_in(wire_d10_41),.data_out(wire_d10_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101043(.data_in(wire_d10_42),.data_out(wire_d10_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101044(.data_in(wire_d10_43),.data_out(wire_d10_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101045(.data_in(wire_d10_44),.data_out(wire_d10_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101046(.data_in(wire_d10_45),.data_out(wire_d10_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101047(.data_in(wire_d10_46),.data_out(wire_d10_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101048(.data_in(wire_d10_47),.data_out(wire_d10_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101049(.data_in(wire_d10_48),.data_out(wire_d10_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101050(.data_in(wire_d10_49),.data_out(wire_d10_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101051(.data_in(wire_d10_50),.data_out(wire_d10_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101052(.data_in(wire_d10_51),.data_out(wire_d10_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101053(.data_in(wire_d10_52),.data_out(wire_d10_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101054(.data_in(wire_d10_53),.data_out(wire_d10_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101055(.data_in(wire_d10_54),.data_out(wire_d10_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101056(.data_in(wire_d10_55),.data_out(wire_d10_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101057(.data_in(wire_d10_56),.data_out(wire_d10_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101058(.data_in(wire_d10_57),.data_out(wire_d10_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101059(.data_in(wire_d10_58),.data_out(wire_d10_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101060(.data_in(wire_d10_59),.data_out(wire_d10_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101061(.data_in(wire_d10_60),.data_out(wire_d10_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101062(.data_in(wire_d10_61),.data_out(wire_d10_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101063(.data_in(wire_d10_62),.data_out(wire_d10_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101064(.data_in(wire_d10_63),.data_out(wire_d10_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101065(.data_in(wire_d10_64),.data_out(wire_d10_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101066(.data_in(wire_d10_65),.data_out(wire_d10_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101067(.data_in(wire_d10_66),.data_out(wire_d10_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101068(.data_in(wire_d10_67),.data_out(wire_d10_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101069(.data_in(wire_d10_68),.data_out(wire_d10_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101070(.data_in(wire_d10_69),.data_out(wire_d10_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101071(.data_in(wire_d10_70),.data_out(wire_d10_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101072(.data_in(wire_d10_71),.data_out(wire_d10_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101073(.data_in(wire_d10_72),.data_out(wire_d10_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101074(.data_in(wire_d10_73),.data_out(wire_d10_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101075(.data_in(wire_d10_74),.data_out(wire_d10_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101076(.data_in(wire_d10_75),.data_out(wire_d10_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101077(.data_in(wire_d10_76),.data_out(wire_d10_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101078(.data_in(wire_d10_77),.data_out(wire_d10_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101079(.data_in(wire_d10_78),.data_out(d_out10),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance120110(.data_in(d_in11),.data_out(wire_d11_0),.clk(clk),.rst(rst));            //channel 12
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance120111(.data_in(wire_d11_0),.data_out(wire_d11_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance120112(.data_in(wire_d11_1),.data_out(wire_d11_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance120113(.data_in(wire_d11_2),.data_out(wire_d11_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance120114(.data_in(wire_d11_3),.data_out(wire_d11_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance120115(.data_in(wire_d11_4),.data_out(wire_d11_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance120116(.data_in(wire_d11_5),.data_out(wire_d11_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance120117(.data_in(wire_d11_6),.data_out(wire_d11_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance120118(.data_in(wire_d11_7),.data_out(wire_d11_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance120119(.data_in(wire_d11_8),.data_out(wire_d11_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201110(.data_in(wire_d11_9),.data_out(wire_d11_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201111(.data_in(wire_d11_10),.data_out(wire_d11_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201112(.data_in(wire_d11_11),.data_out(wire_d11_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201113(.data_in(wire_d11_12),.data_out(wire_d11_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201114(.data_in(wire_d11_13),.data_out(wire_d11_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201115(.data_in(wire_d11_14),.data_out(wire_d11_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201116(.data_in(wire_d11_15),.data_out(wire_d11_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201117(.data_in(wire_d11_16),.data_out(wire_d11_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201118(.data_in(wire_d11_17),.data_out(wire_d11_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201119(.data_in(wire_d11_18),.data_out(wire_d11_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201120(.data_in(wire_d11_19),.data_out(wire_d11_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201121(.data_in(wire_d11_20),.data_out(wire_d11_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201122(.data_in(wire_d11_21),.data_out(wire_d11_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201123(.data_in(wire_d11_22),.data_out(wire_d11_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201124(.data_in(wire_d11_23),.data_out(wire_d11_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201125(.data_in(wire_d11_24),.data_out(wire_d11_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201126(.data_in(wire_d11_25),.data_out(wire_d11_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201127(.data_in(wire_d11_26),.data_out(wire_d11_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201128(.data_in(wire_d11_27),.data_out(wire_d11_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201129(.data_in(wire_d11_28),.data_out(wire_d11_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201130(.data_in(wire_d11_29),.data_out(wire_d11_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201131(.data_in(wire_d11_30),.data_out(wire_d11_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201132(.data_in(wire_d11_31),.data_out(wire_d11_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201133(.data_in(wire_d11_32),.data_out(wire_d11_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201134(.data_in(wire_d11_33),.data_out(wire_d11_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201135(.data_in(wire_d11_34),.data_out(wire_d11_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201136(.data_in(wire_d11_35),.data_out(wire_d11_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201137(.data_in(wire_d11_36),.data_out(wire_d11_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201138(.data_in(wire_d11_37),.data_out(wire_d11_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201139(.data_in(wire_d11_38),.data_out(wire_d11_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201140(.data_in(wire_d11_39),.data_out(wire_d11_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201141(.data_in(wire_d11_40),.data_out(wire_d11_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201142(.data_in(wire_d11_41),.data_out(wire_d11_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201143(.data_in(wire_d11_42),.data_out(wire_d11_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201144(.data_in(wire_d11_43),.data_out(wire_d11_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201145(.data_in(wire_d11_44),.data_out(wire_d11_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201146(.data_in(wire_d11_45),.data_out(wire_d11_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201147(.data_in(wire_d11_46),.data_out(wire_d11_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201148(.data_in(wire_d11_47),.data_out(wire_d11_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201149(.data_in(wire_d11_48),.data_out(wire_d11_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201150(.data_in(wire_d11_49),.data_out(wire_d11_50),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201151(.data_in(wire_d11_50),.data_out(wire_d11_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201152(.data_in(wire_d11_51),.data_out(wire_d11_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201153(.data_in(wire_d11_52),.data_out(wire_d11_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201154(.data_in(wire_d11_53),.data_out(wire_d11_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201155(.data_in(wire_d11_54),.data_out(wire_d11_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201156(.data_in(wire_d11_55),.data_out(wire_d11_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201157(.data_in(wire_d11_56),.data_out(wire_d11_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201158(.data_in(wire_d11_57),.data_out(wire_d11_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201159(.data_in(wire_d11_58),.data_out(wire_d11_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201160(.data_in(wire_d11_59),.data_out(wire_d11_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201161(.data_in(wire_d11_60),.data_out(wire_d11_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201162(.data_in(wire_d11_61),.data_out(wire_d11_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201163(.data_in(wire_d11_62),.data_out(wire_d11_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201164(.data_in(wire_d11_63),.data_out(wire_d11_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201165(.data_in(wire_d11_64),.data_out(wire_d11_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201166(.data_in(wire_d11_65),.data_out(wire_d11_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201167(.data_in(wire_d11_66),.data_out(wire_d11_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201168(.data_in(wire_d11_67),.data_out(wire_d11_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201169(.data_in(wire_d11_68),.data_out(wire_d11_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201170(.data_in(wire_d11_69),.data_out(wire_d11_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201171(.data_in(wire_d11_70),.data_out(wire_d11_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201172(.data_in(wire_d11_71),.data_out(wire_d11_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201173(.data_in(wire_d11_72),.data_out(wire_d11_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201174(.data_in(wire_d11_73),.data_out(wire_d11_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201175(.data_in(wire_d11_74),.data_out(wire_d11_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201176(.data_in(wire_d11_75),.data_out(wire_d11_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201177(.data_in(wire_d11_76),.data_out(wire_d11_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201178(.data_in(wire_d11_77),.data_out(wire_d11_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201179(.data_in(wire_d11_78),.data_out(d_out11),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance130120(.data_in(d_in12),.data_out(wire_d12_0),.clk(clk),.rst(rst));            //channel 13
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance130121(.data_in(wire_d12_0),.data_out(wire_d12_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance130122(.data_in(wire_d12_1),.data_out(wire_d12_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance130123(.data_in(wire_d12_2),.data_out(wire_d12_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance130124(.data_in(wire_d12_3),.data_out(wire_d12_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance130125(.data_in(wire_d12_4),.data_out(wire_d12_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance130126(.data_in(wire_d12_5),.data_out(wire_d12_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance130127(.data_in(wire_d12_6),.data_out(wire_d12_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance130128(.data_in(wire_d12_7),.data_out(wire_d12_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance130129(.data_in(wire_d12_8),.data_out(wire_d12_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301210(.data_in(wire_d12_9),.data_out(wire_d12_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301211(.data_in(wire_d12_10),.data_out(wire_d12_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301212(.data_in(wire_d12_11),.data_out(wire_d12_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301213(.data_in(wire_d12_12),.data_out(wire_d12_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301214(.data_in(wire_d12_13),.data_out(wire_d12_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301215(.data_in(wire_d12_14),.data_out(wire_d12_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301216(.data_in(wire_d12_15),.data_out(wire_d12_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301217(.data_in(wire_d12_16),.data_out(wire_d12_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301218(.data_in(wire_d12_17),.data_out(wire_d12_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301219(.data_in(wire_d12_18),.data_out(wire_d12_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301220(.data_in(wire_d12_19),.data_out(wire_d12_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301221(.data_in(wire_d12_20),.data_out(wire_d12_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301222(.data_in(wire_d12_21),.data_out(wire_d12_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301223(.data_in(wire_d12_22),.data_out(wire_d12_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301224(.data_in(wire_d12_23),.data_out(wire_d12_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301225(.data_in(wire_d12_24),.data_out(wire_d12_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301226(.data_in(wire_d12_25),.data_out(wire_d12_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301227(.data_in(wire_d12_26),.data_out(wire_d12_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301228(.data_in(wire_d12_27),.data_out(wire_d12_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301229(.data_in(wire_d12_28),.data_out(wire_d12_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301230(.data_in(wire_d12_29),.data_out(wire_d12_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301231(.data_in(wire_d12_30),.data_out(wire_d12_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301232(.data_in(wire_d12_31),.data_out(wire_d12_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301233(.data_in(wire_d12_32),.data_out(wire_d12_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301234(.data_in(wire_d12_33),.data_out(wire_d12_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301235(.data_in(wire_d12_34),.data_out(wire_d12_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301236(.data_in(wire_d12_35),.data_out(wire_d12_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301237(.data_in(wire_d12_36),.data_out(wire_d12_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301238(.data_in(wire_d12_37),.data_out(wire_d12_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301239(.data_in(wire_d12_38),.data_out(wire_d12_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301240(.data_in(wire_d12_39),.data_out(wire_d12_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301241(.data_in(wire_d12_40),.data_out(wire_d12_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301242(.data_in(wire_d12_41),.data_out(wire_d12_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301243(.data_in(wire_d12_42),.data_out(wire_d12_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301244(.data_in(wire_d12_43),.data_out(wire_d12_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301245(.data_in(wire_d12_44),.data_out(wire_d12_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301246(.data_in(wire_d12_45),.data_out(wire_d12_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301247(.data_in(wire_d12_46),.data_out(wire_d12_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301248(.data_in(wire_d12_47),.data_out(wire_d12_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301249(.data_in(wire_d12_48),.data_out(wire_d12_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301250(.data_in(wire_d12_49),.data_out(wire_d12_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301251(.data_in(wire_d12_50),.data_out(wire_d12_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301252(.data_in(wire_d12_51),.data_out(wire_d12_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301253(.data_in(wire_d12_52),.data_out(wire_d12_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301254(.data_in(wire_d12_53),.data_out(wire_d12_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301255(.data_in(wire_d12_54),.data_out(wire_d12_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301256(.data_in(wire_d12_55),.data_out(wire_d12_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301257(.data_in(wire_d12_56),.data_out(wire_d12_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301258(.data_in(wire_d12_57),.data_out(wire_d12_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301259(.data_in(wire_d12_58),.data_out(wire_d12_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301260(.data_in(wire_d12_59),.data_out(wire_d12_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301261(.data_in(wire_d12_60),.data_out(wire_d12_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301262(.data_in(wire_d12_61),.data_out(wire_d12_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301263(.data_in(wire_d12_62),.data_out(wire_d12_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301264(.data_in(wire_d12_63),.data_out(wire_d12_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301265(.data_in(wire_d12_64),.data_out(wire_d12_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301266(.data_in(wire_d12_65),.data_out(wire_d12_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301267(.data_in(wire_d12_66),.data_out(wire_d12_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301268(.data_in(wire_d12_67),.data_out(wire_d12_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301269(.data_in(wire_d12_68),.data_out(wire_d12_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301270(.data_in(wire_d12_69),.data_out(wire_d12_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301271(.data_in(wire_d12_70),.data_out(wire_d12_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301272(.data_in(wire_d12_71),.data_out(wire_d12_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301273(.data_in(wire_d12_72),.data_out(wire_d12_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301274(.data_in(wire_d12_73),.data_out(wire_d12_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301275(.data_in(wire_d12_74),.data_out(wire_d12_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301276(.data_in(wire_d12_75),.data_out(wire_d12_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301277(.data_in(wire_d12_76),.data_out(wire_d12_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301278(.data_in(wire_d12_77),.data_out(wire_d12_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301279(.data_in(wire_d12_78),.data_out(d_out12),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance140130(.data_in(d_in13),.data_out(wire_d13_0),.clk(clk),.rst(rst));            //channel 14
	large_adder #(.WIDTH(WIDTH)) large_adder_instance140131(.data_in(wire_d13_0),.data_out(wire_d13_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance140132(.data_in(wire_d13_1),.data_out(wire_d13_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance140133(.data_in(wire_d13_2),.data_out(wire_d13_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance140134(.data_in(wire_d13_3),.data_out(wire_d13_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance140135(.data_in(wire_d13_4),.data_out(wire_d13_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance140136(.data_in(wire_d13_5),.data_out(wire_d13_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance140137(.data_in(wire_d13_6),.data_out(wire_d13_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance140138(.data_in(wire_d13_7),.data_out(wire_d13_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance140139(.data_in(wire_d13_8),.data_out(wire_d13_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401310(.data_in(wire_d13_9),.data_out(wire_d13_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401311(.data_in(wire_d13_10),.data_out(wire_d13_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401312(.data_in(wire_d13_11),.data_out(wire_d13_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401313(.data_in(wire_d13_12),.data_out(wire_d13_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401314(.data_in(wire_d13_13),.data_out(wire_d13_14),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401315(.data_in(wire_d13_14),.data_out(wire_d13_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401316(.data_in(wire_d13_15),.data_out(wire_d13_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401317(.data_in(wire_d13_16),.data_out(wire_d13_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401318(.data_in(wire_d13_17),.data_out(wire_d13_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401319(.data_in(wire_d13_18),.data_out(wire_d13_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401320(.data_in(wire_d13_19),.data_out(wire_d13_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401321(.data_in(wire_d13_20),.data_out(wire_d13_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401322(.data_in(wire_d13_21),.data_out(wire_d13_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401323(.data_in(wire_d13_22),.data_out(wire_d13_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401324(.data_in(wire_d13_23),.data_out(wire_d13_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401325(.data_in(wire_d13_24),.data_out(wire_d13_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401326(.data_in(wire_d13_25),.data_out(wire_d13_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401327(.data_in(wire_d13_26),.data_out(wire_d13_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401328(.data_in(wire_d13_27),.data_out(wire_d13_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401329(.data_in(wire_d13_28),.data_out(wire_d13_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401330(.data_in(wire_d13_29),.data_out(wire_d13_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401331(.data_in(wire_d13_30),.data_out(wire_d13_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401332(.data_in(wire_d13_31),.data_out(wire_d13_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401333(.data_in(wire_d13_32),.data_out(wire_d13_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401334(.data_in(wire_d13_33),.data_out(wire_d13_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401335(.data_in(wire_d13_34),.data_out(wire_d13_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401336(.data_in(wire_d13_35),.data_out(wire_d13_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401337(.data_in(wire_d13_36),.data_out(wire_d13_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401338(.data_in(wire_d13_37),.data_out(wire_d13_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401339(.data_in(wire_d13_38),.data_out(wire_d13_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401340(.data_in(wire_d13_39),.data_out(wire_d13_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401341(.data_in(wire_d13_40),.data_out(wire_d13_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401342(.data_in(wire_d13_41),.data_out(wire_d13_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401343(.data_in(wire_d13_42),.data_out(wire_d13_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401344(.data_in(wire_d13_43),.data_out(wire_d13_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401345(.data_in(wire_d13_44),.data_out(wire_d13_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401346(.data_in(wire_d13_45),.data_out(wire_d13_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401347(.data_in(wire_d13_46),.data_out(wire_d13_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401348(.data_in(wire_d13_47),.data_out(wire_d13_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401349(.data_in(wire_d13_48),.data_out(wire_d13_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401350(.data_in(wire_d13_49),.data_out(wire_d13_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401351(.data_in(wire_d13_50),.data_out(wire_d13_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401352(.data_in(wire_d13_51),.data_out(wire_d13_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401353(.data_in(wire_d13_52),.data_out(wire_d13_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401354(.data_in(wire_d13_53),.data_out(wire_d13_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401355(.data_in(wire_d13_54),.data_out(wire_d13_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401356(.data_in(wire_d13_55),.data_out(wire_d13_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401357(.data_in(wire_d13_56),.data_out(wire_d13_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401358(.data_in(wire_d13_57),.data_out(wire_d13_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401359(.data_in(wire_d13_58),.data_out(wire_d13_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401360(.data_in(wire_d13_59),.data_out(wire_d13_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401361(.data_in(wire_d13_60),.data_out(wire_d13_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401362(.data_in(wire_d13_61),.data_out(wire_d13_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401363(.data_in(wire_d13_62),.data_out(wire_d13_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401364(.data_in(wire_d13_63),.data_out(wire_d13_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401365(.data_in(wire_d13_64),.data_out(wire_d13_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401366(.data_in(wire_d13_65),.data_out(wire_d13_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401367(.data_in(wire_d13_66),.data_out(wire_d13_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401368(.data_in(wire_d13_67),.data_out(wire_d13_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401369(.data_in(wire_d13_68),.data_out(wire_d13_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401370(.data_in(wire_d13_69),.data_out(wire_d13_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401371(.data_in(wire_d13_70),.data_out(wire_d13_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401372(.data_in(wire_d13_71),.data_out(wire_d13_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401373(.data_in(wire_d13_72),.data_out(wire_d13_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401374(.data_in(wire_d13_73),.data_out(wire_d13_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401375(.data_in(wire_d13_74),.data_out(wire_d13_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401376(.data_in(wire_d13_75),.data_out(wire_d13_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401377(.data_in(wire_d13_76),.data_out(wire_d13_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401378(.data_in(wire_d13_77),.data_out(wire_d13_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401379(.data_in(wire_d13_78),.data_out(d_out13),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance150140(.data_in(d_in14),.data_out(wire_d14_0),.clk(clk),.rst(rst));            //channel 15
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance150141(.data_in(wire_d14_0),.data_out(wire_d14_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance150142(.data_in(wire_d14_1),.data_out(wire_d14_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance150143(.data_in(wire_d14_2),.data_out(wire_d14_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance150144(.data_in(wire_d14_3),.data_out(wire_d14_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance150145(.data_in(wire_d14_4),.data_out(wire_d14_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance150146(.data_in(wire_d14_5),.data_out(wire_d14_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance150147(.data_in(wire_d14_6),.data_out(wire_d14_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance150148(.data_in(wire_d14_7),.data_out(wire_d14_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance150149(.data_in(wire_d14_8),.data_out(wire_d14_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501410(.data_in(wire_d14_9),.data_out(wire_d14_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501411(.data_in(wire_d14_10),.data_out(wire_d14_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501412(.data_in(wire_d14_11),.data_out(wire_d14_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501413(.data_in(wire_d14_12),.data_out(wire_d14_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501414(.data_in(wire_d14_13),.data_out(wire_d14_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501415(.data_in(wire_d14_14),.data_out(wire_d14_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501416(.data_in(wire_d14_15),.data_out(wire_d14_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501417(.data_in(wire_d14_16),.data_out(wire_d14_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501418(.data_in(wire_d14_17),.data_out(wire_d14_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501419(.data_in(wire_d14_18),.data_out(wire_d14_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501420(.data_in(wire_d14_19),.data_out(wire_d14_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501421(.data_in(wire_d14_20),.data_out(wire_d14_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501422(.data_in(wire_d14_21),.data_out(wire_d14_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501423(.data_in(wire_d14_22),.data_out(wire_d14_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501424(.data_in(wire_d14_23),.data_out(wire_d14_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501425(.data_in(wire_d14_24),.data_out(wire_d14_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501426(.data_in(wire_d14_25),.data_out(wire_d14_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501427(.data_in(wire_d14_26),.data_out(wire_d14_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501428(.data_in(wire_d14_27),.data_out(wire_d14_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501429(.data_in(wire_d14_28),.data_out(wire_d14_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501430(.data_in(wire_d14_29),.data_out(wire_d14_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501431(.data_in(wire_d14_30),.data_out(wire_d14_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501432(.data_in(wire_d14_31),.data_out(wire_d14_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501433(.data_in(wire_d14_32),.data_out(wire_d14_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501434(.data_in(wire_d14_33),.data_out(wire_d14_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501435(.data_in(wire_d14_34),.data_out(wire_d14_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501436(.data_in(wire_d14_35),.data_out(wire_d14_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501437(.data_in(wire_d14_36),.data_out(wire_d14_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501438(.data_in(wire_d14_37),.data_out(wire_d14_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501439(.data_in(wire_d14_38),.data_out(wire_d14_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501440(.data_in(wire_d14_39),.data_out(wire_d14_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501441(.data_in(wire_d14_40),.data_out(wire_d14_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501442(.data_in(wire_d14_41),.data_out(wire_d14_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501443(.data_in(wire_d14_42),.data_out(wire_d14_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501444(.data_in(wire_d14_43),.data_out(wire_d14_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501445(.data_in(wire_d14_44),.data_out(wire_d14_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501446(.data_in(wire_d14_45),.data_out(wire_d14_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501447(.data_in(wire_d14_46),.data_out(wire_d14_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501448(.data_in(wire_d14_47),.data_out(wire_d14_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501449(.data_in(wire_d14_48),.data_out(wire_d14_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501450(.data_in(wire_d14_49),.data_out(wire_d14_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501451(.data_in(wire_d14_50),.data_out(wire_d14_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501452(.data_in(wire_d14_51),.data_out(wire_d14_52),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501453(.data_in(wire_d14_52),.data_out(wire_d14_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501454(.data_in(wire_d14_53),.data_out(wire_d14_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501455(.data_in(wire_d14_54),.data_out(wire_d14_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501456(.data_in(wire_d14_55),.data_out(wire_d14_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501457(.data_in(wire_d14_56),.data_out(wire_d14_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501458(.data_in(wire_d14_57),.data_out(wire_d14_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501459(.data_in(wire_d14_58),.data_out(wire_d14_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501460(.data_in(wire_d14_59),.data_out(wire_d14_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501461(.data_in(wire_d14_60),.data_out(wire_d14_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501462(.data_in(wire_d14_61),.data_out(wire_d14_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501463(.data_in(wire_d14_62),.data_out(wire_d14_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501464(.data_in(wire_d14_63),.data_out(wire_d14_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501465(.data_in(wire_d14_64),.data_out(wire_d14_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501466(.data_in(wire_d14_65),.data_out(wire_d14_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501467(.data_in(wire_d14_66),.data_out(wire_d14_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501468(.data_in(wire_d14_67),.data_out(wire_d14_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501469(.data_in(wire_d14_68),.data_out(wire_d14_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501470(.data_in(wire_d14_69),.data_out(wire_d14_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501471(.data_in(wire_d14_70),.data_out(wire_d14_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501472(.data_in(wire_d14_71),.data_out(wire_d14_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501473(.data_in(wire_d14_72),.data_out(wire_d14_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501474(.data_in(wire_d14_73),.data_out(wire_d14_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501475(.data_in(wire_d14_74),.data_out(wire_d14_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501476(.data_in(wire_d14_75),.data_out(wire_d14_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501477(.data_in(wire_d14_76),.data_out(wire_d14_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501478(.data_in(wire_d14_77),.data_out(wire_d14_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501479(.data_in(wire_d14_78),.data_out(d_out14),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance160150(.data_in(d_in15),.data_out(wire_d15_0),.clk(clk),.rst(rst));            //channel 16
	register #(.WIDTH(WIDTH)) register_instance160151(.data_in(wire_d15_0),.data_out(wire_d15_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance160152(.data_in(wire_d15_1),.data_out(wire_d15_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance160153(.data_in(wire_d15_2),.data_out(wire_d15_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance160154(.data_in(wire_d15_3),.data_out(wire_d15_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance160155(.data_in(wire_d15_4),.data_out(wire_d15_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance160156(.data_in(wire_d15_5),.data_out(wire_d15_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance160157(.data_in(wire_d15_6),.data_out(wire_d15_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance160158(.data_in(wire_d15_7),.data_out(wire_d15_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance160159(.data_in(wire_d15_8),.data_out(wire_d15_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601510(.data_in(wire_d15_9),.data_out(wire_d15_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601511(.data_in(wire_d15_10),.data_out(wire_d15_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601512(.data_in(wire_d15_11),.data_out(wire_d15_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601513(.data_in(wire_d15_12),.data_out(wire_d15_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601514(.data_in(wire_d15_13),.data_out(wire_d15_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601515(.data_in(wire_d15_14),.data_out(wire_d15_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601516(.data_in(wire_d15_15),.data_out(wire_d15_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601517(.data_in(wire_d15_16),.data_out(wire_d15_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601518(.data_in(wire_d15_17),.data_out(wire_d15_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601519(.data_in(wire_d15_18),.data_out(wire_d15_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601520(.data_in(wire_d15_19),.data_out(wire_d15_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601521(.data_in(wire_d15_20),.data_out(wire_d15_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601522(.data_in(wire_d15_21),.data_out(wire_d15_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601523(.data_in(wire_d15_22),.data_out(wire_d15_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601524(.data_in(wire_d15_23),.data_out(wire_d15_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601525(.data_in(wire_d15_24),.data_out(wire_d15_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601526(.data_in(wire_d15_25),.data_out(wire_d15_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601527(.data_in(wire_d15_26),.data_out(wire_d15_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601528(.data_in(wire_d15_27),.data_out(wire_d15_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601529(.data_in(wire_d15_28),.data_out(wire_d15_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601530(.data_in(wire_d15_29),.data_out(wire_d15_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601531(.data_in(wire_d15_30),.data_out(wire_d15_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601532(.data_in(wire_d15_31),.data_out(wire_d15_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601533(.data_in(wire_d15_32),.data_out(wire_d15_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601534(.data_in(wire_d15_33),.data_out(wire_d15_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601535(.data_in(wire_d15_34),.data_out(wire_d15_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601536(.data_in(wire_d15_35),.data_out(wire_d15_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601537(.data_in(wire_d15_36),.data_out(wire_d15_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601538(.data_in(wire_d15_37),.data_out(wire_d15_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601539(.data_in(wire_d15_38),.data_out(wire_d15_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601540(.data_in(wire_d15_39),.data_out(wire_d15_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601541(.data_in(wire_d15_40),.data_out(wire_d15_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601542(.data_in(wire_d15_41),.data_out(wire_d15_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601543(.data_in(wire_d15_42),.data_out(wire_d15_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601544(.data_in(wire_d15_43),.data_out(wire_d15_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601545(.data_in(wire_d15_44),.data_out(wire_d15_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601546(.data_in(wire_d15_45),.data_out(wire_d15_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601547(.data_in(wire_d15_46),.data_out(wire_d15_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601548(.data_in(wire_d15_47),.data_out(wire_d15_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601549(.data_in(wire_d15_48),.data_out(wire_d15_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601550(.data_in(wire_d15_49),.data_out(wire_d15_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601551(.data_in(wire_d15_50),.data_out(wire_d15_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601552(.data_in(wire_d15_51),.data_out(wire_d15_52),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601553(.data_in(wire_d15_52),.data_out(wire_d15_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601554(.data_in(wire_d15_53),.data_out(wire_d15_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601555(.data_in(wire_d15_54),.data_out(wire_d15_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601556(.data_in(wire_d15_55),.data_out(wire_d15_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601557(.data_in(wire_d15_56),.data_out(wire_d15_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601558(.data_in(wire_d15_57),.data_out(wire_d15_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601559(.data_in(wire_d15_58),.data_out(wire_d15_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601560(.data_in(wire_d15_59),.data_out(wire_d15_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601561(.data_in(wire_d15_60),.data_out(wire_d15_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601562(.data_in(wire_d15_61),.data_out(wire_d15_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601563(.data_in(wire_d15_62),.data_out(wire_d15_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601564(.data_in(wire_d15_63),.data_out(wire_d15_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601565(.data_in(wire_d15_64),.data_out(wire_d15_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601566(.data_in(wire_d15_65),.data_out(wire_d15_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601567(.data_in(wire_d15_66),.data_out(wire_d15_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601568(.data_in(wire_d15_67),.data_out(wire_d15_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601569(.data_in(wire_d15_68),.data_out(wire_d15_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601570(.data_in(wire_d15_69),.data_out(wire_d15_70),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601571(.data_in(wire_d15_70),.data_out(wire_d15_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601572(.data_in(wire_d15_71),.data_out(wire_d15_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601573(.data_in(wire_d15_72),.data_out(wire_d15_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601574(.data_in(wire_d15_73),.data_out(wire_d15_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601575(.data_in(wire_d15_74),.data_out(wire_d15_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601576(.data_in(wire_d15_75),.data_out(wire_d15_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601577(.data_in(wire_d15_76),.data_out(wire_d15_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601578(.data_in(wire_d15_77),.data_out(wire_d15_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601579(.data_in(wire_d15_78),.data_out(d_out15),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance170160(.data_in(d_in16),.data_out(wire_d16_0),.clk(clk),.rst(rst));            //channel 17
	large_mux #(.WIDTH(WIDTH)) large_mux_instance170161(.data_in(wire_d16_0),.data_out(wire_d16_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance170162(.data_in(wire_d16_1),.data_out(wire_d16_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance170163(.data_in(wire_d16_2),.data_out(wire_d16_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance170164(.data_in(wire_d16_3),.data_out(wire_d16_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance170165(.data_in(wire_d16_4),.data_out(wire_d16_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance170166(.data_in(wire_d16_5),.data_out(wire_d16_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance170167(.data_in(wire_d16_6),.data_out(wire_d16_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance170168(.data_in(wire_d16_7),.data_out(wire_d16_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance170169(.data_in(wire_d16_8),.data_out(wire_d16_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701610(.data_in(wire_d16_9),.data_out(wire_d16_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701611(.data_in(wire_d16_10),.data_out(wire_d16_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701612(.data_in(wire_d16_11),.data_out(wire_d16_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701613(.data_in(wire_d16_12),.data_out(wire_d16_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701614(.data_in(wire_d16_13),.data_out(wire_d16_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701615(.data_in(wire_d16_14),.data_out(wire_d16_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701616(.data_in(wire_d16_15),.data_out(wire_d16_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701617(.data_in(wire_d16_16),.data_out(wire_d16_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701618(.data_in(wire_d16_17),.data_out(wire_d16_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701619(.data_in(wire_d16_18),.data_out(wire_d16_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701620(.data_in(wire_d16_19),.data_out(wire_d16_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701621(.data_in(wire_d16_20),.data_out(wire_d16_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701622(.data_in(wire_d16_21),.data_out(wire_d16_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701623(.data_in(wire_d16_22),.data_out(wire_d16_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701624(.data_in(wire_d16_23),.data_out(wire_d16_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701625(.data_in(wire_d16_24),.data_out(wire_d16_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701626(.data_in(wire_d16_25),.data_out(wire_d16_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701627(.data_in(wire_d16_26),.data_out(wire_d16_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701628(.data_in(wire_d16_27),.data_out(wire_d16_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701629(.data_in(wire_d16_28),.data_out(wire_d16_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701630(.data_in(wire_d16_29),.data_out(wire_d16_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701631(.data_in(wire_d16_30),.data_out(wire_d16_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701632(.data_in(wire_d16_31),.data_out(wire_d16_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701633(.data_in(wire_d16_32),.data_out(wire_d16_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701634(.data_in(wire_d16_33),.data_out(wire_d16_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701635(.data_in(wire_d16_34),.data_out(wire_d16_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701636(.data_in(wire_d16_35),.data_out(wire_d16_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701637(.data_in(wire_d16_36),.data_out(wire_d16_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701638(.data_in(wire_d16_37),.data_out(wire_d16_38),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701639(.data_in(wire_d16_38),.data_out(wire_d16_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701640(.data_in(wire_d16_39),.data_out(wire_d16_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701641(.data_in(wire_d16_40),.data_out(wire_d16_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701642(.data_in(wire_d16_41),.data_out(wire_d16_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701643(.data_in(wire_d16_42),.data_out(wire_d16_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701644(.data_in(wire_d16_43),.data_out(wire_d16_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701645(.data_in(wire_d16_44),.data_out(wire_d16_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701646(.data_in(wire_d16_45),.data_out(wire_d16_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701647(.data_in(wire_d16_46),.data_out(wire_d16_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701648(.data_in(wire_d16_47),.data_out(wire_d16_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701649(.data_in(wire_d16_48),.data_out(wire_d16_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701650(.data_in(wire_d16_49),.data_out(wire_d16_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701651(.data_in(wire_d16_50),.data_out(wire_d16_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701652(.data_in(wire_d16_51),.data_out(wire_d16_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701653(.data_in(wire_d16_52),.data_out(wire_d16_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701654(.data_in(wire_d16_53),.data_out(wire_d16_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701655(.data_in(wire_d16_54),.data_out(wire_d16_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701656(.data_in(wire_d16_55),.data_out(wire_d16_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701657(.data_in(wire_d16_56),.data_out(wire_d16_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701658(.data_in(wire_d16_57),.data_out(wire_d16_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701659(.data_in(wire_d16_58),.data_out(wire_d16_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701660(.data_in(wire_d16_59),.data_out(wire_d16_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701661(.data_in(wire_d16_60),.data_out(wire_d16_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701662(.data_in(wire_d16_61),.data_out(wire_d16_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701663(.data_in(wire_d16_62),.data_out(wire_d16_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701664(.data_in(wire_d16_63),.data_out(wire_d16_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701665(.data_in(wire_d16_64),.data_out(wire_d16_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701666(.data_in(wire_d16_65),.data_out(wire_d16_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701667(.data_in(wire_d16_66),.data_out(wire_d16_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701668(.data_in(wire_d16_67),.data_out(wire_d16_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701669(.data_in(wire_d16_68),.data_out(wire_d16_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701670(.data_in(wire_d16_69),.data_out(wire_d16_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701671(.data_in(wire_d16_70),.data_out(wire_d16_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701672(.data_in(wire_d16_71),.data_out(wire_d16_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701673(.data_in(wire_d16_72),.data_out(wire_d16_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701674(.data_in(wire_d16_73),.data_out(wire_d16_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701675(.data_in(wire_d16_74),.data_out(wire_d16_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701676(.data_in(wire_d16_75),.data_out(wire_d16_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701677(.data_in(wire_d16_76),.data_out(wire_d16_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701678(.data_in(wire_d16_77),.data_out(wire_d16_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701679(.data_in(wire_d16_78),.data_out(d_out16),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance180170(.data_in(d_in17),.data_out(wire_d17_0),.clk(clk),.rst(rst));            //channel 18
	encoder #(.WIDTH(WIDTH)) encoder_instance180171(.data_in(wire_d17_0),.data_out(wire_d17_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance180172(.data_in(wire_d17_1),.data_out(wire_d17_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance180173(.data_in(wire_d17_2),.data_out(wire_d17_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance180174(.data_in(wire_d17_3),.data_out(wire_d17_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance180175(.data_in(wire_d17_4),.data_out(wire_d17_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance180176(.data_in(wire_d17_5),.data_out(wire_d17_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance180177(.data_in(wire_d17_6),.data_out(wire_d17_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance180178(.data_in(wire_d17_7),.data_out(wire_d17_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance180179(.data_in(wire_d17_8),.data_out(wire_d17_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801710(.data_in(wire_d17_9),.data_out(wire_d17_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801711(.data_in(wire_d17_10),.data_out(wire_d17_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801712(.data_in(wire_d17_11),.data_out(wire_d17_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801713(.data_in(wire_d17_12),.data_out(wire_d17_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801714(.data_in(wire_d17_13),.data_out(wire_d17_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801715(.data_in(wire_d17_14),.data_out(wire_d17_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801716(.data_in(wire_d17_15),.data_out(wire_d17_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801717(.data_in(wire_d17_16),.data_out(wire_d17_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801718(.data_in(wire_d17_17),.data_out(wire_d17_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801719(.data_in(wire_d17_18),.data_out(wire_d17_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801720(.data_in(wire_d17_19),.data_out(wire_d17_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801721(.data_in(wire_d17_20),.data_out(wire_d17_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801722(.data_in(wire_d17_21),.data_out(wire_d17_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801723(.data_in(wire_d17_22),.data_out(wire_d17_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801724(.data_in(wire_d17_23),.data_out(wire_d17_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801725(.data_in(wire_d17_24),.data_out(wire_d17_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801726(.data_in(wire_d17_25),.data_out(wire_d17_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801727(.data_in(wire_d17_26),.data_out(wire_d17_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801728(.data_in(wire_d17_27),.data_out(wire_d17_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801729(.data_in(wire_d17_28),.data_out(wire_d17_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801730(.data_in(wire_d17_29),.data_out(wire_d17_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801731(.data_in(wire_d17_30),.data_out(wire_d17_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801732(.data_in(wire_d17_31),.data_out(wire_d17_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801733(.data_in(wire_d17_32),.data_out(wire_d17_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801734(.data_in(wire_d17_33),.data_out(wire_d17_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801735(.data_in(wire_d17_34),.data_out(wire_d17_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801736(.data_in(wire_d17_35),.data_out(wire_d17_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801737(.data_in(wire_d17_36),.data_out(wire_d17_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801738(.data_in(wire_d17_37),.data_out(wire_d17_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801739(.data_in(wire_d17_38),.data_out(wire_d17_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801740(.data_in(wire_d17_39),.data_out(wire_d17_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801741(.data_in(wire_d17_40),.data_out(wire_d17_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801742(.data_in(wire_d17_41),.data_out(wire_d17_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801743(.data_in(wire_d17_42),.data_out(wire_d17_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801744(.data_in(wire_d17_43),.data_out(wire_d17_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801745(.data_in(wire_d17_44),.data_out(wire_d17_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801746(.data_in(wire_d17_45),.data_out(wire_d17_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801747(.data_in(wire_d17_46),.data_out(wire_d17_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801748(.data_in(wire_d17_47),.data_out(wire_d17_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801749(.data_in(wire_d17_48),.data_out(wire_d17_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801750(.data_in(wire_d17_49),.data_out(wire_d17_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801751(.data_in(wire_d17_50),.data_out(wire_d17_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801752(.data_in(wire_d17_51),.data_out(wire_d17_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801753(.data_in(wire_d17_52),.data_out(wire_d17_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801754(.data_in(wire_d17_53),.data_out(wire_d17_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801755(.data_in(wire_d17_54),.data_out(wire_d17_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801756(.data_in(wire_d17_55),.data_out(wire_d17_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801757(.data_in(wire_d17_56),.data_out(wire_d17_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801758(.data_in(wire_d17_57),.data_out(wire_d17_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801759(.data_in(wire_d17_58),.data_out(wire_d17_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801760(.data_in(wire_d17_59),.data_out(wire_d17_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801761(.data_in(wire_d17_60),.data_out(wire_d17_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801762(.data_in(wire_d17_61),.data_out(wire_d17_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801763(.data_in(wire_d17_62),.data_out(wire_d17_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801764(.data_in(wire_d17_63),.data_out(wire_d17_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801765(.data_in(wire_d17_64),.data_out(wire_d17_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801766(.data_in(wire_d17_65),.data_out(wire_d17_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801767(.data_in(wire_d17_66),.data_out(wire_d17_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801768(.data_in(wire_d17_67),.data_out(wire_d17_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801769(.data_in(wire_d17_68),.data_out(wire_d17_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801770(.data_in(wire_d17_69),.data_out(wire_d17_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801771(.data_in(wire_d17_70),.data_out(wire_d17_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801772(.data_in(wire_d17_71),.data_out(wire_d17_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801773(.data_in(wire_d17_72),.data_out(wire_d17_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801774(.data_in(wire_d17_73),.data_out(wire_d17_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801775(.data_in(wire_d17_74),.data_out(wire_d17_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801776(.data_in(wire_d17_75),.data_out(wire_d17_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801777(.data_in(wire_d17_76),.data_out(wire_d17_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801778(.data_in(wire_d17_77),.data_out(wire_d17_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801779(.data_in(wire_d17_78),.data_out(d_out17),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance190180(.data_in(d_in18),.data_out(wire_d18_0),.clk(clk),.rst(rst));            //channel 19
	large_adder #(.WIDTH(WIDTH)) large_adder_instance190181(.data_in(wire_d18_0),.data_out(wire_d18_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance190182(.data_in(wire_d18_1),.data_out(wire_d18_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance190183(.data_in(wire_d18_2),.data_out(wire_d18_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance190184(.data_in(wire_d18_3),.data_out(wire_d18_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance190185(.data_in(wire_d18_4),.data_out(wire_d18_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance190186(.data_in(wire_d18_5),.data_out(wire_d18_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance190187(.data_in(wire_d18_6),.data_out(wire_d18_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance190188(.data_in(wire_d18_7),.data_out(wire_d18_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance190189(.data_in(wire_d18_8),.data_out(wire_d18_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901810(.data_in(wire_d18_9),.data_out(wire_d18_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901811(.data_in(wire_d18_10),.data_out(wire_d18_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901812(.data_in(wire_d18_11),.data_out(wire_d18_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901813(.data_in(wire_d18_12),.data_out(wire_d18_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901814(.data_in(wire_d18_13),.data_out(wire_d18_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901815(.data_in(wire_d18_14),.data_out(wire_d18_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901816(.data_in(wire_d18_15),.data_out(wire_d18_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901817(.data_in(wire_d18_16),.data_out(wire_d18_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901818(.data_in(wire_d18_17),.data_out(wire_d18_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901819(.data_in(wire_d18_18),.data_out(wire_d18_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901820(.data_in(wire_d18_19),.data_out(wire_d18_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901821(.data_in(wire_d18_20),.data_out(wire_d18_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901822(.data_in(wire_d18_21),.data_out(wire_d18_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901823(.data_in(wire_d18_22),.data_out(wire_d18_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901824(.data_in(wire_d18_23),.data_out(wire_d18_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901825(.data_in(wire_d18_24),.data_out(wire_d18_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901826(.data_in(wire_d18_25),.data_out(wire_d18_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901827(.data_in(wire_d18_26),.data_out(wire_d18_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901828(.data_in(wire_d18_27),.data_out(wire_d18_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901829(.data_in(wire_d18_28),.data_out(wire_d18_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901830(.data_in(wire_d18_29),.data_out(wire_d18_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901831(.data_in(wire_d18_30),.data_out(wire_d18_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901832(.data_in(wire_d18_31),.data_out(wire_d18_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901833(.data_in(wire_d18_32),.data_out(wire_d18_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901834(.data_in(wire_d18_33),.data_out(wire_d18_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901835(.data_in(wire_d18_34),.data_out(wire_d18_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901836(.data_in(wire_d18_35),.data_out(wire_d18_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901837(.data_in(wire_d18_36),.data_out(wire_d18_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901838(.data_in(wire_d18_37),.data_out(wire_d18_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901839(.data_in(wire_d18_38),.data_out(wire_d18_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901840(.data_in(wire_d18_39),.data_out(wire_d18_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901841(.data_in(wire_d18_40),.data_out(wire_d18_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901842(.data_in(wire_d18_41),.data_out(wire_d18_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901843(.data_in(wire_d18_42),.data_out(wire_d18_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901844(.data_in(wire_d18_43),.data_out(wire_d18_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901845(.data_in(wire_d18_44),.data_out(wire_d18_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901846(.data_in(wire_d18_45),.data_out(wire_d18_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901847(.data_in(wire_d18_46),.data_out(wire_d18_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901848(.data_in(wire_d18_47),.data_out(wire_d18_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901849(.data_in(wire_d18_48),.data_out(wire_d18_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901850(.data_in(wire_d18_49),.data_out(wire_d18_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901851(.data_in(wire_d18_50),.data_out(wire_d18_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901852(.data_in(wire_d18_51),.data_out(wire_d18_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901853(.data_in(wire_d18_52),.data_out(wire_d18_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901854(.data_in(wire_d18_53),.data_out(wire_d18_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901855(.data_in(wire_d18_54),.data_out(wire_d18_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901856(.data_in(wire_d18_55),.data_out(wire_d18_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901857(.data_in(wire_d18_56),.data_out(wire_d18_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901858(.data_in(wire_d18_57),.data_out(wire_d18_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901859(.data_in(wire_d18_58),.data_out(wire_d18_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901860(.data_in(wire_d18_59),.data_out(wire_d18_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901861(.data_in(wire_d18_60),.data_out(wire_d18_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901862(.data_in(wire_d18_61),.data_out(wire_d18_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901863(.data_in(wire_d18_62),.data_out(wire_d18_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901864(.data_in(wire_d18_63),.data_out(wire_d18_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901865(.data_in(wire_d18_64),.data_out(wire_d18_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901866(.data_in(wire_d18_65),.data_out(wire_d18_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901867(.data_in(wire_d18_66),.data_out(wire_d18_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901868(.data_in(wire_d18_67),.data_out(wire_d18_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901869(.data_in(wire_d18_68),.data_out(wire_d18_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901870(.data_in(wire_d18_69),.data_out(wire_d18_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901871(.data_in(wire_d18_70),.data_out(wire_d18_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901872(.data_in(wire_d18_71),.data_out(wire_d18_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901873(.data_in(wire_d18_72),.data_out(wire_d18_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901874(.data_in(wire_d18_73),.data_out(wire_d18_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901875(.data_in(wire_d18_74),.data_out(wire_d18_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901876(.data_in(wire_d18_75),.data_out(wire_d18_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901877(.data_in(wire_d18_76),.data_out(wire_d18_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901878(.data_in(wire_d18_77),.data_out(wire_d18_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901879(.data_in(wire_d18_78),.data_out(d_out18),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance200190(.data_in(d_in19),.data_out(wire_d19_0),.clk(clk),.rst(rst));            //channel 20
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance200191(.data_in(wire_d19_0),.data_out(wire_d19_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance200192(.data_in(wire_d19_1),.data_out(wire_d19_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance200193(.data_in(wire_d19_2),.data_out(wire_d19_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance200194(.data_in(wire_d19_3),.data_out(wire_d19_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance200195(.data_in(wire_d19_4),.data_out(wire_d19_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance200196(.data_in(wire_d19_5),.data_out(wire_d19_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance200197(.data_in(wire_d19_6),.data_out(wire_d19_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance200198(.data_in(wire_d19_7),.data_out(wire_d19_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance200199(.data_in(wire_d19_8),.data_out(wire_d19_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001910(.data_in(wire_d19_9),.data_out(wire_d19_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001911(.data_in(wire_d19_10),.data_out(wire_d19_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001912(.data_in(wire_d19_11),.data_out(wire_d19_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001913(.data_in(wire_d19_12),.data_out(wire_d19_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001914(.data_in(wire_d19_13),.data_out(wire_d19_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001915(.data_in(wire_d19_14),.data_out(wire_d19_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001916(.data_in(wire_d19_15),.data_out(wire_d19_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001917(.data_in(wire_d19_16),.data_out(wire_d19_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001918(.data_in(wire_d19_17),.data_out(wire_d19_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001919(.data_in(wire_d19_18),.data_out(wire_d19_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001920(.data_in(wire_d19_19),.data_out(wire_d19_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001921(.data_in(wire_d19_20),.data_out(wire_d19_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001922(.data_in(wire_d19_21),.data_out(wire_d19_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001923(.data_in(wire_d19_22),.data_out(wire_d19_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001924(.data_in(wire_d19_23),.data_out(wire_d19_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001925(.data_in(wire_d19_24),.data_out(wire_d19_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001926(.data_in(wire_d19_25),.data_out(wire_d19_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001927(.data_in(wire_d19_26),.data_out(wire_d19_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001928(.data_in(wire_d19_27),.data_out(wire_d19_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001929(.data_in(wire_d19_28),.data_out(wire_d19_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001930(.data_in(wire_d19_29),.data_out(wire_d19_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001931(.data_in(wire_d19_30),.data_out(wire_d19_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001932(.data_in(wire_d19_31),.data_out(wire_d19_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001933(.data_in(wire_d19_32),.data_out(wire_d19_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001934(.data_in(wire_d19_33),.data_out(wire_d19_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001935(.data_in(wire_d19_34),.data_out(wire_d19_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001936(.data_in(wire_d19_35),.data_out(wire_d19_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001937(.data_in(wire_d19_36),.data_out(wire_d19_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001938(.data_in(wire_d19_37),.data_out(wire_d19_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001939(.data_in(wire_d19_38),.data_out(wire_d19_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001940(.data_in(wire_d19_39),.data_out(wire_d19_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001941(.data_in(wire_d19_40),.data_out(wire_d19_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001942(.data_in(wire_d19_41),.data_out(wire_d19_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001943(.data_in(wire_d19_42),.data_out(wire_d19_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001944(.data_in(wire_d19_43),.data_out(wire_d19_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001945(.data_in(wire_d19_44),.data_out(wire_d19_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001946(.data_in(wire_d19_45),.data_out(wire_d19_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001947(.data_in(wire_d19_46),.data_out(wire_d19_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001948(.data_in(wire_d19_47),.data_out(wire_d19_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001949(.data_in(wire_d19_48),.data_out(wire_d19_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001950(.data_in(wire_d19_49),.data_out(wire_d19_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001951(.data_in(wire_d19_50),.data_out(wire_d19_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001952(.data_in(wire_d19_51),.data_out(wire_d19_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001953(.data_in(wire_d19_52),.data_out(wire_d19_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001954(.data_in(wire_d19_53),.data_out(wire_d19_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001955(.data_in(wire_d19_54),.data_out(wire_d19_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001956(.data_in(wire_d19_55),.data_out(wire_d19_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001957(.data_in(wire_d19_56),.data_out(wire_d19_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001958(.data_in(wire_d19_57),.data_out(wire_d19_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001959(.data_in(wire_d19_58),.data_out(wire_d19_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001960(.data_in(wire_d19_59),.data_out(wire_d19_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001961(.data_in(wire_d19_60),.data_out(wire_d19_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001962(.data_in(wire_d19_61),.data_out(wire_d19_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001963(.data_in(wire_d19_62),.data_out(wire_d19_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001964(.data_in(wire_d19_63),.data_out(wire_d19_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001965(.data_in(wire_d19_64),.data_out(wire_d19_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001966(.data_in(wire_d19_65),.data_out(wire_d19_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001967(.data_in(wire_d19_66),.data_out(wire_d19_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001968(.data_in(wire_d19_67),.data_out(wire_d19_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001969(.data_in(wire_d19_68),.data_out(wire_d19_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001970(.data_in(wire_d19_69),.data_out(wire_d19_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001971(.data_in(wire_d19_70),.data_out(wire_d19_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001972(.data_in(wire_d19_71),.data_out(wire_d19_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001973(.data_in(wire_d19_72),.data_out(wire_d19_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001974(.data_in(wire_d19_73),.data_out(wire_d19_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001975(.data_in(wire_d19_74),.data_out(wire_d19_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001976(.data_in(wire_d19_75),.data_out(wire_d19_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001977(.data_in(wire_d19_76),.data_out(wire_d19_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001978(.data_in(wire_d19_77),.data_out(wire_d19_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001979(.data_in(wire_d19_78),.data_out(d_out19),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance210200(.data_in(d_in20),.data_out(wire_d20_0),.clk(clk),.rst(rst));            //channel 21
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance210201(.data_in(wire_d20_0),.data_out(wire_d20_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance210202(.data_in(wire_d20_1),.data_out(wire_d20_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance210203(.data_in(wire_d20_2),.data_out(wire_d20_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance210204(.data_in(wire_d20_3),.data_out(wire_d20_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance210205(.data_in(wire_d20_4),.data_out(wire_d20_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance210206(.data_in(wire_d20_5),.data_out(wire_d20_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance210207(.data_in(wire_d20_6),.data_out(wire_d20_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance210208(.data_in(wire_d20_7),.data_out(wire_d20_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance210209(.data_in(wire_d20_8),.data_out(wire_d20_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102010(.data_in(wire_d20_9),.data_out(wire_d20_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102011(.data_in(wire_d20_10),.data_out(wire_d20_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102012(.data_in(wire_d20_11),.data_out(wire_d20_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102013(.data_in(wire_d20_12),.data_out(wire_d20_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102014(.data_in(wire_d20_13),.data_out(wire_d20_14),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102015(.data_in(wire_d20_14),.data_out(wire_d20_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102016(.data_in(wire_d20_15),.data_out(wire_d20_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102017(.data_in(wire_d20_16),.data_out(wire_d20_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102018(.data_in(wire_d20_17),.data_out(wire_d20_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102019(.data_in(wire_d20_18),.data_out(wire_d20_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102020(.data_in(wire_d20_19),.data_out(wire_d20_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102021(.data_in(wire_d20_20),.data_out(wire_d20_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102022(.data_in(wire_d20_21),.data_out(wire_d20_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102023(.data_in(wire_d20_22),.data_out(wire_d20_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102024(.data_in(wire_d20_23),.data_out(wire_d20_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102025(.data_in(wire_d20_24),.data_out(wire_d20_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102026(.data_in(wire_d20_25),.data_out(wire_d20_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102027(.data_in(wire_d20_26),.data_out(wire_d20_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102028(.data_in(wire_d20_27),.data_out(wire_d20_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102029(.data_in(wire_d20_28),.data_out(wire_d20_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102030(.data_in(wire_d20_29),.data_out(wire_d20_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102031(.data_in(wire_d20_30),.data_out(wire_d20_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102032(.data_in(wire_d20_31),.data_out(wire_d20_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102033(.data_in(wire_d20_32),.data_out(wire_d20_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102034(.data_in(wire_d20_33),.data_out(wire_d20_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102035(.data_in(wire_d20_34),.data_out(wire_d20_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102036(.data_in(wire_d20_35),.data_out(wire_d20_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102037(.data_in(wire_d20_36),.data_out(wire_d20_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102038(.data_in(wire_d20_37),.data_out(wire_d20_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102039(.data_in(wire_d20_38),.data_out(wire_d20_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102040(.data_in(wire_d20_39),.data_out(wire_d20_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102041(.data_in(wire_d20_40),.data_out(wire_d20_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102042(.data_in(wire_d20_41),.data_out(wire_d20_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102043(.data_in(wire_d20_42),.data_out(wire_d20_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102044(.data_in(wire_d20_43),.data_out(wire_d20_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102045(.data_in(wire_d20_44),.data_out(wire_d20_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102046(.data_in(wire_d20_45),.data_out(wire_d20_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102047(.data_in(wire_d20_46),.data_out(wire_d20_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102048(.data_in(wire_d20_47),.data_out(wire_d20_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102049(.data_in(wire_d20_48),.data_out(wire_d20_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102050(.data_in(wire_d20_49),.data_out(wire_d20_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102051(.data_in(wire_d20_50),.data_out(wire_d20_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102052(.data_in(wire_d20_51),.data_out(wire_d20_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102053(.data_in(wire_d20_52),.data_out(wire_d20_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102054(.data_in(wire_d20_53),.data_out(wire_d20_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102055(.data_in(wire_d20_54),.data_out(wire_d20_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102056(.data_in(wire_d20_55),.data_out(wire_d20_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102057(.data_in(wire_d20_56),.data_out(wire_d20_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102058(.data_in(wire_d20_57),.data_out(wire_d20_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102059(.data_in(wire_d20_58),.data_out(wire_d20_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102060(.data_in(wire_d20_59),.data_out(wire_d20_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102061(.data_in(wire_d20_60),.data_out(wire_d20_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102062(.data_in(wire_d20_61),.data_out(wire_d20_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102063(.data_in(wire_d20_62),.data_out(wire_d20_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102064(.data_in(wire_d20_63),.data_out(wire_d20_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102065(.data_in(wire_d20_64),.data_out(wire_d20_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102066(.data_in(wire_d20_65),.data_out(wire_d20_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102067(.data_in(wire_d20_66),.data_out(wire_d20_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102068(.data_in(wire_d20_67),.data_out(wire_d20_68),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102069(.data_in(wire_d20_68),.data_out(wire_d20_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102070(.data_in(wire_d20_69),.data_out(wire_d20_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102071(.data_in(wire_d20_70),.data_out(wire_d20_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102072(.data_in(wire_d20_71),.data_out(wire_d20_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102073(.data_in(wire_d20_72),.data_out(wire_d20_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102074(.data_in(wire_d20_73),.data_out(wire_d20_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102075(.data_in(wire_d20_74),.data_out(wire_d20_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102076(.data_in(wire_d20_75),.data_out(wire_d20_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102077(.data_in(wire_d20_76),.data_out(wire_d20_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102078(.data_in(wire_d20_77),.data_out(wire_d20_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102079(.data_in(wire_d20_78),.data_out(d_out20),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance220210(.data_in(d_in21),.data_out(wire_d21_0),.clk(clk),.rst(rst));            //channel 22
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance220211(.data_in(wire_d21_0),.data_out(wire_d21_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance220212(.data_in(wire_d21_1),.data_out(wire_d21_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance220213(.data_in(wire_d21_2),.data_out(wire_d21_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance220214(.data_in(wire_d21_3),.data_out(wire_d21_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance220215(.data_in(wire_d21_4),.data_out(wire_d21_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance220216(.data_in(wire_d21_5),.data_out(wire_d21_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance220217(.data_in(wire_d21_6),.data_out(wire_d21_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance220218(.data_in(wire_d21_7),.data_out(wire_d21_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance220219(.data_in(wire_d21_8),.data_out(wire_d21_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202110(.data_in(wire_d21_9),.data_out(wire_d21_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202111(.data_in(wire_d21_10),.data_out(wire_d21_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202112(.data_in(wire_d21_11),.data_out(wire_d21_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202113(.data_in(wire_d21_12),.data_out(wire_d21_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202114(.data_in(wire_d21_13),.data_out(wire_d21_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202115(.data_in(wire_d21_14),.data_out(wire_d21_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202116(.data_in(wire_d21_15),.data_out(wire_d21_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202117(.data_in(wire_d21_16),.data_out(wire_d21_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202118(.data_in(wire_d21_17),.data_out(wire_d21_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202119(.data_in(wire_d21_18),.data_out(wire_d21_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202120(.data_in(wire_d21_19),.data_out(wire_d21_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202121(.data_in(wire_d21_20),.data_out(wire_d21_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202122(.data_in(wire_d21_21),.data_out(wire_d21_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202123(.data_in(wire_d21_22),.data_out(wire_d21_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202124(.data_in(wire_d21_23),.data_out(wire_d21_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202125(.data_in(wire_d21_24),.data_out(wire_d21_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202126(.data_in(wire_d21_25),.data_out(wire_d21_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202127(.data_in(wire_d21_26),.data_out(wire_d21_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202128(.data_in(wire_d21_27),.data_out(wire_d21_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202129(.data_in(wire_d21_28),.data_out(wire_d21_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202130(.data_in(wire_d21_29),.data_out(wire_d21_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202131(.data_in(wire_d21_30),.data_out(wire_d21_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202132(.data_in(wire_d21_31),.data_out(wire_d21_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202133(.data_in(wire_d21_32),.data_out(wire_d21_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202134(.data_in(wire_d21_33),.data_out(wire_d21_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202135(.data_in(wire_d21_34),.data_out(wire_d21_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202136(.data_in(wire_d21_35),.data_out(wire_d21_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202137(.data_in(wire_d21_36),.data_out(wire_d21_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202138(.data_in(wire_d21_37),.data_out(wire_d21_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202139(.data_in(wire_d21_38),.data_out(wire_d21_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202140(.data_in(wire_d21_39),.data_out(wire_d21_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202141(.data_in(wire_d21_40),.data_out(wire_d21_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202142(.data_in(wire_d21_41),.data_out(wire_d21_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202143(.data_in(wire_d21_42),.data_out(wire_d21_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202144(.data_in(wire_d21_43),.data_out(wire_d21_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202145(.data_in(wire_d21_44),.data_out(wire_d21_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202146(.data_in(wire_d21_45),.data_out(wire_d21_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202147(.data_in(wire_d21_46),.data_out(wire_d21_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202148(.data_in(wire_d21_47),.data_out(wire_d21_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202149(.data_in(wire_d21_48),.data_out(wire_d21_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202150(.data_in(wire_d21_49),.data_out(wire_d21_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202151(.data_in(wire_d21_50),.data_out(wire_d21_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202152(.data_in(wire_d21_51),.data_out(wire_d21_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202153(.data_in(wire_d21_52),.data_out(wire_d21_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202154(.data_in(wire_d21_53),.data_out(wire_d21_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202155(.data_in(wire_d21_54),.data_out(wire_d21_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202156(.data_in(wire_d21_55),.data_out(wire_d21_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202157(.data_in(wire_d21_56),.data_out(wire_d21_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202158(.data_in(wire_d21_57),.data_out(wire_d21_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202159(.data_in(wire_d21_58),.data_out(wire_d21_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202160(.data_in(wire_d21_59),.data_out(wire_d21_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202161(.data_in(wire_d21_60),.data_out(wire_d21_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202162(.data_in(wire_d21_61),.data_out(wire_d21_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202163(.data_in(wire_d21_62),.data_out(wire_d21_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202164(.data_in(wire_d21_63),.data_out(wire_d21_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202165(.data_in(wire_d21_64),.data_out(wire_d21_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202166(.data_in(wire_d21_65),.data_out(wire_d21_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202167(.data_in(wire_d21_66),.data_out(wire_d21_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202168(.data_in(wire_d21_67),.data_out(wire_d21_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202169(.data_in(wire_d21_68),.data_out(wire_d21_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202170(.data_in(wire_d21_69),.data_out(wire_d21_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202171(.data_in(wire_d21_70),.data_out(wire_d21_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202172(.data_in(wire_d21_71),.data_out(wire_d21_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202173(.data_in(wire_d21_72),.data_out(wire_d21_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202174(.data_in(wire_d21_73),.data_out(wire_d21_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202175(.data_in(wire_d21_74),.data_out(wire_d21_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202176(.data_in(wire_d21_75),.data_out(wire_d21_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202177(.data_in(wire_d21_76),.data_out(wire_d21_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202178(.data_in(wire_d21_77),.data_out(wire_d21_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202179(.data_in(wire_d21_78),.data_out(d_out21),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance230220(.data_in(d_in22),.data_out(wire_d22_0),.clk(clk),.rst(rst));            //channel 23
	large_mux #(.WIDTH(WIDTH)) large_mux_instance230221(.data_in(wire_d22_0),.data_out(wire_d22_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance230222(.data_in(wire_d22_1),.data_out(wire_d22_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance230223(.data_in(wire_d22_2),.data_out(wire_d22_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance230224(.data_in(wire_d22_3),.data_out(wire_d22_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance230225(.data_in(wire_d22_4),.data_out(wire_d22_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance230226(.data_in(wire_d22_5),.data_out(wire_d22_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance230227(.data_in(wire_d22_6),.data_out(wire_d22_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance230228(.data_in(wire_d22_7),.data_out(wire_d22_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance230229(.data_in(wire_d22_8),.data_out(wire_d22_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302210(.data_in(wire_d22_9),.data_out(wire_d22_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302211(.data_in(wire_d22_10),.data_out(wire_d22_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302212(.data_in(wire_d22_11),.data_out(wire_d22_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302213(.data_in(wire_d22_12),.data_out(wire_d22_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302214(.data_in(wire_d22_13),.data_out(wire_d22_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302215(.data_in(wire_d22_14),.data_out(wire_d22_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302216(.data_in(wire_d22_15),.data_out(wire_d22_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302217(.data_in(wire_d22_16),.data_out(wire_d22_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302218(.data_in(wire_d22_17),.data_out(wire_d22_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302219(.data_in(wire_d22_18),.data_out(wire_d22_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302220(.data_in(wire_d22_19),.data_out(wire_d22_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302221(.data_in(wire_d22_20),.data_out(wire_d22_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302222(.data_in(wire_d22_21),.data_out(wire_d22_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302223(.data_in(wire_d22_22),.data_out(wire_d22_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302224(.data_in(wire_d22_23),.data_out(wire_d22_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302225(.data_in(wire_d22_24),.data_out(wire_d22_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302226(.data_in(wire_d22_25),.data_out(wire_d22_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302227(.data_in(wire_d22_26),.data_out(wire_d22_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302228(.data_in(wire_d22_27),.data_out(wire_d22_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302229(.data_in(wire_d22_28),.data_out(wire_d22_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302230(.data_in(wire_d22_29),.data_out(wire_d22_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302231(.data_in(wire_d22_30),.data_out(wire_d22_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302232(.data_in(wire_d22_31),.data_out(wire_d22_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302233(.data_in(wire_d22_32),.data_out(wire_d22_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302234(.data_in(wire_d22_33),.data_out(wire_d22_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302235(.data_in(wire_d22_34),.data_out(wire_d22_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302236(.data_in(wire_d22_35),.data_out(wire_d22_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302237(.data_in(wire_d22_36),.data_out(wire_d22_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302238(.data_in(wire_d22_37),.data_out(wire_d22_38),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302239(.data_in(wire_d22_38),.data_out(wire_d22_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302240(.data_in(wire_d22_39),.data_out(wire_d22_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302241(.data_in(wire_d22_40),.data_out(wire_d22_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302242(.data_in(wire_d22_41),.data_out(wire_d22_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302243(.data_in(wire_d22_42),.data_out(wire_d22_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302244(.data_in(wire_d22_43),.data_out(wire_d22_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302245(.data_in(wire_d22_44),.data_out(wire_d22_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302246(.data_in(wire_d22_45),.data_out(wire_d22_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302247(.data_in(wire_d22_46),.data_out(wire_d22_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302248(.data_in(wire_d22_47),.data_out(wire_d22_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302249(.data_in(wire_d22_48),.data_out(wire_d22_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302250(.data_in(wire_d22_49),.data_out(wire_d22_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302251(.data_in(wire_d22_50),.data_out(wire_d22_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302252(.data_in(wire_d22_51),.data_out(wire_d22_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302253(.data_in(wire_d22_52),.data_out(wire_d22_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302254(.data_in(wire_d22_53),.data_out(wire_d22_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302255(.data_in(wire_d22_54),.data_out(wire_d22_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302256(.data_in(wire_d22_55),.data_out(wire_d22_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302257(.data_in(wire_d22_56),.data_out(wire_d22_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302258(.data_in(wire_d22_57),.data_out(wire_d22_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302259(.data_in(wire_d22_58),.data_out(wire_d22_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302260(.data_in(wire_d22_59),.data_out(wire_d22_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302261(.data_in(wire_d22_60),.data_out(wire_d22_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302262(.data_in(wire_d22_61),.data_out(wire_d22_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302263(.data_in(wire_d22_62),.data_out(wire_d22_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302264(.data_in(wire_d22_63),.data_out(wire_d22_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302265(.data_in(wire_d22_64),.data_out(wire_d22_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302266(.data_in(wire_d22_65),.data_out(wire_d22_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302267(.data_in(wire_d22_66),.data_out(wire_d22_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302268(.data_in(wire_d22_67),.data_out(wire_d22_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302269(.data_in(wire_d22_68),.data_out(wire_d22_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302270(.data_in(wire_d22_69),.data_out(wire_d22_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302271(.data_in(wire_d22_70),.data_out(wire_d22_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302272(.data_in(wire_d22_71),.data_out(wire_d22_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302273(.data_in(wire_d22_72),.data_out(wire_d22_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302274(.data_in(wire_d22_73),.data_out(wire_d22_74),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302275(.data_in(wire_d22_74),.data_out(wire_d22_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302276(.data_in(wire_d22_75),.data_out(wire_d22_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302277(.data_in(wire_d22_76),.data_out(wire_d22_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302278(.data_in(wire_d22_77),.data_out(wire_d22_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302279(.data_in(wire_d22_78),.data_out(d_out22),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance240230(.data_in(d_in23),.data_out(wire_d23_0),.clk(clk),.rst(rst));            //channel 24
	register #(.WIDTH(WIDTH)) register_instance240231(.data_in(wire_d23_0),.data_out(wire_d23_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance240232(.data_in(wire_d23_1),.data_out(wire_d23_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance240233(.data_in(wire_d23_2),.data_out(wire_d23_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance240234(.data_in(wire_d23_3),.data_out(wire_d23_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance240235(.data_in(wire_d23_4),.data_out(wire_d23_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance240236(.data_in(wire_d23_5),.data_out(wire_d23_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance240237(.data_in(wire_d23_6),.data_out(wire_d23_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance240238(.data_in(wire_d23_7),.data_out(wire_d23_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance240239(.data_in(wire_d23_8),.data_out(wire_d23_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402310(.data_in(wire_d23_9),.data_out(wire_d23_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402311(.data_in(wire_d23_10),.data_out(wire_d23_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402312(.data_in(wire_d23_11),.data_out(wire_d23_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402313(.data_in(wire_d23_12),.data_out(wire_d23_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402314(.data_in(wire_d23_13),.data_out(wire_d23_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402315(.data_in(wire_d23_14),.data_out(wire_d23_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402316(.data_in(wire_d23_15),.data_out(wire_d23_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402317(.data_in(wire_d23_16),.data_out(wire_d23_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402318(.data_in(wire_d23_17),.data_out(wire_d23_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402319(.data_in(wire_d23_18),.data_out(wire_d23_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402320(.data_in(wire_d23_19),.data_out(wire_d23_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402321(.data_in(wire_d23_20),.data_out(wire_d23_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402322(.data_in(wire_d23_21),.data_out(wire_d23_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402323(.data_in(wire_d23_22),.data_out(wire_d23_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402324(.data_in(wire_d23_23),.data_out(wire_d23_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402325(.data_in(wire_d23_24),.data_out(wire_d23_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402326(.data_in(wire_d23_25),.data_out(wire_d23_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402327(.data_in(wire_d23_26),.data_out(wire_d23_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402328(.data_in(wire_d23_27),.data_out(wire_d23_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402329(.data_in(wire_d23_28),.data_out(wire_d23_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402330(.data_in(wire_d23_29),.data_out(wire_d23_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402331(.data_in(wire_d23_30),.data_out(wire_d23_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402332(.data_in(wire_d23_31),.data_out(wire_d23_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402333(.data_in(wire_d23_32),.data_out(wire_d23_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402334(.data_in(wire_d23_33),.data_out(wire_d23_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402335(.data_in(wire_d23_34),.data_out(wire_d23_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402336(.data_in(wire_d23_35),.data_out(wire_d23_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402337(.data_in(wire_d23_36),.data_out(wire_d23_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402338(.data_in(wire_d23_37),.data_out(wire_d23_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402339(.data_in(wire_d23_38),.data_out(wire_d23_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402340(.data_in(wire_d23_39),.data_out(wire_d23_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402341(.data_in(wire_d23_40),.data_out(wire_d23_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402342(.data_in(wire_d23_41),.data_out(wire_d23_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402343(.data_in(wire_d23_42),.data_out(wire_d23_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402344(.data_in(wire_d23_43),.data_out(wire_d23_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402345(.data_in(wire_d23_44),.data_out(wire_d23_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402346(.data_in(wire_d23_45),.data_out(wire_d23_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402347(.data_in(wire_d23_46),.data_out(wire_d23_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402348(.data_in(wire_d23_47),.data_out(wire_d23_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402349(.data_in(wire_d23_48),.data_out(wire_d23_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402350(.data_in(wire_d23_49),.data_out(wire_d23_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402351(.data_in(wire_d23_50),.data_out(wire_d23_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402352(.data_in(wire_d23_51),.data_out(wire_d23_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402353(.data_in(wire_d23_52),.data_out(wire_d23_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402354(.data_in(wire_d23_53),.data_out(wire_d23_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402355(.data_in(wire_d23_54),.data_out(wire_d23_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402356(.data_in(wire_d23_55),.data_out(wire_d23_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402357(.data_in(wire_d23_56),.data_out(wire_d23_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402358(.data_in(wire_d23_57),.data_out(wire_d23_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402359(.data_in(wire_d23_58),.data_out(wire_d23_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402360(.data_in(wire_d23_59),.data_out(wire_d23_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402361(.data_in(wire_d23_60),.data_out(wire_d23_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402362(.data_in(wire_d23_61),.data_out(wire_d23_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402363(.data_in(wire_d23_62),.data_out(wire_d23_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402364(.data_in(wire_d23_63),.data_out(wire_d23_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402365(.data_in(wire_d23_64),.data_out(wire_d23_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402366(.data_in(wire_d23_65),.data_out(wire_d23_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402367(.data_in(wire_d23_66),.data_out(wire_d23_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402368(.data_in(wire_d23_67),.data_out(wire_d23_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402369(.data_in(wire_d23_68),.data_out(wire_d23_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402370(.data_in(wire_d23_69),.data_out(wire_d23_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402371(.data_in(wire_d23_70),.data_out(wire_d23_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402372(.data_in(wire_d23_71),.data_out(wire_d23_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402373(.data_in(wire_d23_72),.data_out(wire_d23_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402374(.data_in(wire_d23_73),.data_out(wire_d23_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402375(.data_in(wire_d23_74),.data_out(wire_d23_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402376(.data_in(wire_d23_75),.data_out(wire_d23_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402377(.data_in(wire_d23_76),.data_out(wire_d23_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402378(.data_in(wire_d23_77),.data_out(wire_d23_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402379(.data_in(wire_d23_78),.data_out(d_out23),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance250240(.data_in(d_in24),.data_out(wire_d24_0),.clk(clk),.rst(rst));            //channel 25
	large_mux #(.WIDTH(WIDTH)) large_mux_instance250241(.data_in(wire_d24_0),.data_out(wire_d24_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance250242(.data_in(wire_d24_1),.data_out(wire_d24_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance250243(.data_in(wire_d24_2),.data_out(wire_d24_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance250244(.data_in(wire_d24_3),.data_out(wire_d24_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance250245(.data_in(wire_d24_4),.data_out(wire_d24_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance250246(.data_in(wire_d24_5),.data_out(wire_d24_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance250247(.data_in(wire_d24_6),.data_out(wire_d24_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance250248(.data_in(wire_d24_7),.data_out(wire_d24_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance250249(.data_in(wire_d24_8),.data_out(wire_d24_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502410(.data_in(wire_d24_9),.data_out(wire_d24_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502411(.data_in(wire_d24_10),.data_out(wire_d24_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502412(.data_in(wire_d24_11),.data_out(wire_d24_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502413(.data_in(wire_d24_12),.data_out(wire_d24_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502414(.data_in(wire_d24_13),.data_out(wire_d24_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502415(.data_in(wire_d24_14),.data_out(wire_d24_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502416(.data_in(wire_d24_15),.data_out(wire_d24_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502417(.data_in(wire_d24_16),.data_out(wire_d24_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502418(.data_in(wire_d24_17),.data_out(wire_d24_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502419(.data_in(wire_d24_18),.data_out(wire_d24_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502420(.data_in(wire_d24_19),.data_out(wire_d24_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502421(.data_in(wire_d24_20),.data_out(wire_d24_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502422(.data_in(wire_d24_21),.data_out(wire_d24_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502423(.data_in(wire_d24_22),.data_out(wire_d24_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502424(.data_in(wire_d24_23),.data_out(wire_d24_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502425(.data_in(wire_d24_24),.data_out(wire_d24_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502426(.data_in(wire_d24_25),.data_out(wire_d24_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502427(.data_in(wire_d24_26),.data_out(wire_d24_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502428(.data_in(wire_d24_27),.data_out(wire_d24_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502429(.data_in(wire_d24_28),.data_out(wire_d24_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502430(.data_in(wire_d24_29),.data_out(wire_d24_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502431(.data_in(wire_d24_30),.data_out(wire_d24_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502432(.data_in(wire_d24_31),.data_out(wire_d24_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502433(.data_in(wire_d24_32),.data_out(wire_d24_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502434(.data_in(wire_d24_33),.data_out(wire_d24_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502435(.data_in(wire_d24_34),.data_out(wire_d24_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502436(.data_in(wire_d24_35),.data_out(wire_d24_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502437(.data_in(wire_d24_36),.data_out(wire_d24_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502438(.data_in(wire_d24_37),.data_out(wire_d24_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502439(.data_in(wire_d24_38),.data_out(wire_d24_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502440(.data_in(wire_d24_39),.data_out(wire_d24_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502441(.data_in(wire_d24_40),.data_out(wire_d24_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502442(.data_in(wire_d24_41),.data_out(wire_d24_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502443(.data_in(wire_d24_42),.data_out(wire_d24_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502444(.data_in(wire_d24_43),.data_out(wire_d24_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502445(.data_in(wire_d24_44),.data_out(wire_d24_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502446(.data_in(wire_d24_45),.data_out(wire_d24_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502447(.data_in(wire_d24_46),.data_out(wire_d24_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502448(.data_in(wire_d24_47),.data_out(wire_d24_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502449(.data_in(wire_d24_48),.data_out(wire_d24_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502450(.data_in(wire_d24_49),.data_out(wire_d24_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502451(.data_in(wire_d24_50),.data_out(wire_d24_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502452(.data_in(wire_d24_51),.data_out(wire_d24_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502453(.data_in(wire_d24_52),.data_out(wire_d24_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502454(.data_in(wire_d24_53),.data_out(wire_d24_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502455(.data_in(wire_d24_54),.data_out(wire_d24_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502456(.data_in(wire_d24_55),.data_out(wire_d24_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502457(.data_in(wire_d24_56),.data_out(wire_d24_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502458(.data_in(wire_d24_57),.data_out(wire_d24_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502459(.data_in(wire_d24_58),.data_out(wire_d24_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502460(.data_in(wire_d24_59),.data_out(wire_d24_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502461(.data_in(wire_d24_60),.data_out(wire_d24_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502462(.data_in(wire_d24_61),.data_out(wire_d24_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502463(.data_in(wire_d24_62),.data_out(wire_d24_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502464(.data_in(wire_d24_63),.data_out(wire_d24_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502465(.data_in(wire_d24_64),.data_out(wire_d24_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502466(.data_in(wire_d24_65),.data_out(wire_d24_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502467(.data_in(wire_d24_66),.data_out(wire_d24_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502468(.data_in(wire_d24_67),.data_out(wire_d24_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502469(.data_in(wire_d24_68),.data_out(wire_d24_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502470(.data_in(wire_d24_69),.data_out(wire_d24_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502471(.data_in(wire_d24_70),.data_out(wire_d24_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502472(.data_in(wire_d24_71),.data_out(wire_d24_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502473(.data_in(wire_d24_72),.data_out(wire_d24_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502474(.data_in(wire_d24_73),.data_out(wire_d24_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502475(.data_in(wire_d24_74),.data_out(wire_d24_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502476(.data_in(wire_d24_75),.data_out(wire_d24_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502477(.data_in(wire_d24_76),.data_out(wire_d24_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502478(.data_in(wire_d24_77),.data_out(wire_d24_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502479(.data_in(wire_d24_78),.data_out(d_out24),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance260250(.data_in(d_in25),.data_out(wire_d25_0),.clk(clk),.rst(rst));            //channel 26
	encoder #(.WIDTH(WIDTH)) encoder_instance260251(.data_in(wire_d25_0),.data_out(wire_d25_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance260252(.data_in(wire_d25_1),.data_out(wire_d25_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance260253(.data_in(wire_d25_2),.data_out(wire_d25_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance260254(.data_in(wire_d25_3),.data_out(wire_d25_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance260255(.data_in(wire_d25_4),.data_out(wire_d25_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance260256(.data_in(wire_d25_5),.data_out(wire_d25_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance260257(.data_in(wire_d25_6),.data_out(wire_d25_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance260258(.data_in(wire_d25_7),.data_out(wire_d25_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance260259(.data_in(wire_d25_8),.data_out(wire_d25_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602510(.data_in(wire_d25_9),.data_out(wire_d25_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602511(.data_in(wire_d25_10),.data_out(wire_d25_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602512(.data_in(wire_d25_11),.data_out(wire_d25_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602513(.data_in(wire_d25_12),.data_out(wire_d25_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602514(.data_in(wire_d25_13),.data_out(wire_d25_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602515(.data_in(wire_d25_14),.data_out(wire_d25_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602516(.data_in(wire_d25_15),.data_out(wire_d25_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602517(.data_in(wire_d25_16),.data_out(wire_d25_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602518(.data_in(wire_d25_17),.data_out(wire_d25_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602519(.data_in(wire_d25_18),.data_out(wire_d25_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602520(.data_in(wire_d25_19),.data_out(wire_d25_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602521(.data_in(wire_d25_20),.data_out(wire_d25_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602522(.data_in(wire_d25_21),.data_out(wire_d25_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602523(.data_in(wire_d25_22),.data_out(wire_d25_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602524(.data_in(wire_d25_23),.data_out(wire_d25_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602525(.data_in(wire_d25_24),.data_out(wire_d25_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602526(.data_in(wire_d25_25),.data_out(wire_d25_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602527(.data_in(wire_d25_26),.data_out(wire_d25_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602528(.data_in(wire_d25_27),.data_out(wire_d25_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602529(.data_in(wire_d25_28),.data_out(wire_d25_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602530(.data_in(wire_d25_29),.data_out(wire_d25_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602531(.data_in(wire_d25_30),.data_out(wire_d25_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602532(.data_in(wire_d25_31),.data_out(wire_d25_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602533(.data_in(wire_d25_32),.data_out(wire_d25_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602534(.data_in(wire_d25_33),.data_out(wire_d25_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602535(.data_in(wire_d25_34),.data_out(wire_d25_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602536(.data_in(wire_d25_35),.data_out(wire_d25_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602537(.data_in(wire_d25_36),.data_out(wire_d25_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602538(.data_in(wire_d25_37),.data_out(wire_d25_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602539(.data_in(wire_d25_38),.data_out(wire_d25_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602540(.data_in(wire_d25_39),.data_out(wire_d25_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602541(.data_in(wire_d25_40),.data_out(wire_d25_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602542(.data_in(wire_d25_41),.data_out(wire_d25_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602543(.data_in(wire_d25_42),.data_out(wire_d25_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602544(.data_in(wire_d25_43),.data_out(wire_d25_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602545(.data_in(wire_d25_44),.data_out(wire_d25_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602546(.data_in(wire_d25_45),.data_out(wire_d25_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602547(.data_in(wire_d25_46),.data_out(wire_d25_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602548(.data_in(wire_d25_47),.data_out(wire_d25_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602549(.data_in(wire_d25_48),.data_out(wire_d25_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602550(.data_in(wire_d25_49),.data_out(wire_d25_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602551(.data_in(wire_d25_50),.data_out(wire_d25_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602552(.data_in(wire_d25_51),.data_out(wire_d25_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602553(.data_in(wire_d25_52),.data_out(wire_d25_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602554(.data_in(wire_d25_53),.data_out(wire_d25_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602555(.data_in(wire_d25_54),.data_out(wire_d25_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602556(.data_in(wire_d25_55),.data_out(wire_d25_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602557(.data_in(wire_d25_56),.data_out(wire_d25_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602558(.data_in(wire_d25_57),.data_out(wire_d25_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602559(.data_in(wire_d25_58),.data_out(wire_d25_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602560(.data_in(wire_d25_59),.data_out(wire_d25_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602561(.data_in(wire_d25_60),.data_out(wire_d25_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602562(.data_in(wire_d25_61),.data_out(wire_d25_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602563(.data_in(wire_d25_62),.data_out(wire_d25_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602564(.data_in(wire_d25_63),.data_out(wire_d25_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602565(.data_in(wire_d25_64),.data_out(wire_d25_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602566(.data_in(wire_d25_65),.data_out(wire_d25_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602567(.data_in(wire_d25_66),.data_out(wire_d25_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602568(.data_in(wire_d25_67),.data_out(wire_d25_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602569(.data_in(wire_d25_68),.data_out(wire_d25_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602570(.data_in(wire_d25_69),.data_out(wire_d25_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602571(.data_in(wire_d25_70),.data_out(wire_d25_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602572(.data_in(wire_d25_71),.data_out(wire_d25_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602573(.data_in(wire_d25_72),.data_out(wire_d25_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602574(.data_in(wire_d25_73),.data_out(wire_d25_74),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602575(.data_in(wire_d25_74),.data_out(wire_d25_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602576(.data_in(wire_d25_75),.data_out(wire_d25_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602577(.data_in(wire_d25_76),.data_out(wire_d25_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602578(.data_in(wire_d25_77),.data_out(wire_d25_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602579(.data_in(wire_d25_78),.data_out(d_out25),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance270260(.data_in(d_in26),.data_out(wire_d26_0),.clk(clk),.rst(rst));            //channel 27
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance270261(.data_in(wire_d26_0),.data_out(wire_d26_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance270262(.data_in(wire_d26_1),.data_out(wire_d26_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance270263(.data_in(wire_d26_2),.data_out(wire_d26_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance270264(.data_in(wire_d26_3),.data_out(wire_d26_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance270265(.data_in(wire_d26_4),.data_out(wire_d26_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance270266(.data_in(wire_d26_5),.data_out(wire_d26_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance270267(.data_in(wire_d26_6),.data_out(wire_d26_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance270268(.data_in(wire_d26_7),.data_out(wire_d26_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance270269(.data_in(wire_d26_8),.data_out(wire_d26_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702610(.data_in(wire_d26_9),.data_out(wire_d26_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702611(.data_in(wire_d26_10),.data_out(wire_d26_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702612(.data_in(wire_d26_11),.data_out(wire_d26_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702613(.data_in(wire_d26_12),.data_out(wire_d26_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702614(.data_in(wire_d26_13),.data_out(wire_d26_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702615(.data_in(wire_d26_14),.data_out(wire_d26_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702616(.data_in(wire_d26_15),.data_out(wire_d26_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702617(.data_in(wire_d26_16),.data_out(wire_d26_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702618(.data_in(wire_d26_17),.data_out(wire_d26_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702619(.data_in(wire_d26_18),.data_out(wire_d26_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702620(.data_in(wire_d26_19),.data_out(wire_d26_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702621(.data_in(wire_d26_20),.data_out(wire_d26_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702622(.data_in(wire_d26_21),.data_out(wire_d26_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702623(.data_in(wire_d26_22),.data_out(wire_d26_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702624(.data_in(wire_d26_23),.data_out(wire_d26_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702625(.data_in(wire_d26_24),.data_out(wire_d26_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702626(.data_in(wire_d26_25),.data_out(wire_d26_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702627(.data_in(wire_d26_26),.data_out(wire_d26_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702628(.data_in(wire_d26_27),.data_out(wire_d26_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702629(.data_in(wire_d26_28),.data_out(wire_d26_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702630(.data_in(wire_d26_29),.data_out(wire_d26_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702631(.data_in(wire_d26_30),.data_out(wire_d26_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702632(.data_in(wire_d26_31),.data_out(wire_d26_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702633(.data_in(wire_d26_32),.data_out(wire_d26_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702634(.data_in(wire_d26_33),.data_out(wire_d26_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702635(.data_in(wire_d26_34),.data_out(wire_d26_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702636(.data_in(wire_d26_35),.data_out(wire_d26_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702637(.data_in(wire_d26_36),.data_out(wire_d26_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702638(.data_in(wire_d26_37),.data_out(wire_d26_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702639(.data_in(wire_d26_38),.data_out(wire_d26_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702640(.data_in(wire_d26_39),.data_out(wire_d26_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702641(.data_in(wire_d26_40),.data_out(wire_d26_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702642(.data_in(wire_d26_41),.data_out(wire_d26_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702643(.data_in(wire_d26_42),.data_out(wire_d26_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702644(.data_in(wire_d26_43),.data_out(wire_d26_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702645(.data_in(wire_d26_44),.data_out(wire_d26_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702646(.data_in(wire_d26_45),.data_out(wire_d26_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702647(.data_in(wire_d26_46),.data_out(wire_d26_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702648(.data_in(wire_d26_47),.data_out(wire_d26_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702649(.data_in(wire_d26_48),.data_out(wire_d26_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702650(.data_in(wire_d26_49),.data_out(wire_d26_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702651(.data_in(wire_d26_50),.data_out(wire_d26_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702652(.data_in(wire_d26_51),.data_out(wire_d26_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702653(.data_in(wire_d26_52),.data_out(wire_d26_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702654(.data_in(wire_d26_53),.data_out(wire_d26_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702655(.data_in(wire_d26_54),.data_out(wire_d26_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702656(.data_in(wire_d26_55),.data_out(wire_d26_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702657(.data_in(wire_d26_56),.data_out(wire_d26_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702658(.data_in(wire_d26_57),.data_out(wire_d26_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702659(.data_in(wire_d26_58),.data_out(wire_d26_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702660(.data_in(wire_d26_59),.data_out(wire_d26_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702661(.data_in(wire_d26_60),.data_out(wire_d26_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702662(.data_in(wire_d26_61),.data_out(wire_d26_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702663(.data_in(wire_d26_62),.data_out(wire_d26_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702664(.data_in(wire_d26_63),.data_out(wire_d26_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702665(.data_in(wire_d26_64),.data_out(wire_d26_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702666(.data_in(wire_d26_65),.data_out(wire_d26_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702667(.data_in(wire_d26_66),.data_out(wire_d26_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702668(.data_in(wire_d26_67),.data_out(wire_d26_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702669(.data_in(wire_d26_68),.data_out(wire_d26_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702670(.data_in(wire_d26_69),.data_out(wire_d26_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702671(.data_in(wire_d26_70),.data_out(wire_d26_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702672(.data_in(wire_d26_71),.data_out(wire_d26_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702673(.data_in(wire_d26_72),.data_out(wire_d26_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702674(.data_in(wire_d26_73),.data_out(wire_d26_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702675(.data_in(wire_d26_74),.data_out(wire_d26_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702676(.data_in(wire_d26_75),.data_out(wire_d26_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702677(.data_in(wire_d26_76),.data_out(wire_d26_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702678(.data_in(wire_d26_77),.data_out(wire_d26_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702679(.data_in(wire_d26_78),.data_out(d_out26),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance280270(.data_in(d_in27),.data_out(wire_d27_0),.clk(clk),.rst(rst));            //channel 28
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance280271(.data_in(wire_d27_0),.data_out(wire_d27_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance280272(.data_in(wire_d27_1),.data_out(wire_d27_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance280273(.data_in(wire_d27_2),.data_out(wire_d27_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance280274(.data_in(wire_d27_3),.data_out(wire_d27_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance280275(.data_in(wire_d27_4),.data_out(wire_d27_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance280276(.data_in(wire_d27_5),.data_out(wire_d27_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance280277(.data_in(wire_d27_6),.data_out(wire_d27_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance280278(.data_in(wire_d27_7),.data_out(wire_d27_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance280279(.data_in(wire_d27_8),.data_out(wire_d27_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802710(.data_in(wire_d27_9),.data_out(wire_d27_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802711(.data_in(wire_d27_10),.data_out(wire_d27_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802712(.data_in(wire_d27_11),.data_out(wire_d27_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802713(.data_in(wire_d27_12),.data_out(wire_d27_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802714(.data_in(wire_d27_13),.data_out(wire_d27_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802715(.data_in(wire_d27_14),.data_out(wire_d27_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802716(.data_in(wire_d27_15),.data_out(wire_d27_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802717(.data_in(wire_d27_16),.data_out(wire_d27_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802718(.data_in(wire_d27_17),.data_out(wire_d27_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802719(.data_in(wire_d27_18),.data_out(wire_d27_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802720(.data_in(wire_d27_19),.data_out(wire_d27_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802721(.data_in(wire_d27_20),.data_out(wire_d27_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802722(.data_in(wire_d27_21),.data_out(wire_d27_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802723(.data_in(wire_d27_22),.data_out(wire_d27_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802724(.data_in(wire_d27_23),.data_out(wire_d27_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802725(.data_in(wire_d27_24),.data_out(wire_d27_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802726(.data_in(wire_d27_25),.data_out(wire_d27_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802727(.data_in(wire_d27_26),.data_out(wire_d27_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802728(.data_in(wire_d27_27),.data_out(wire_d27_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802729(.data_in(wire_d27_28),.data_out(wire_d27_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802730(.data_in(wire_d27_29),.data_out(wire_d27_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802731(.data_in(wire_d27_30),.data_out(wire_d27_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802732(.data_in(wire_d27_31),.data_out(wire_d27_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802733(.data_in(wire_d27_32),.data_out(wire_d27_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802734(.data_in(wire_d27_33),.data_out(wire_d27_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802735(.data_in(wire_d27_34),.data_out(wire_d27_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802736(.data_in(wire_d27_35),.data_out(wire_d27_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802737(.data_in(wire_d27_36),.data_out(wire_d27_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802738(.data_in(wire_d27_37),.data_out(wire_d27_38),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802739(.data_in(wire_d27_38),.data_out(wire_d27_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802740(.data_in(wire_d27_39),.data_out(wire_d27_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802741(.data_in(wire_d27_40),.data_out(wire_d27_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802742(.data_in(wire_d27_41),.data_out(wire_d27_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802743(.data_in(wire_d27_42),.data_out(wire_d27_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802744(.data_in(wire_d27_43),.data_out(wire_d27_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802745(.data_in(wire_d27_44),.data_out(wire_d27_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802746(.data_in(wire_d27_45),.data_out(wire_d27_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802747(.data_in(wire_d27_46),.data_out(wire_d27_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802748(.data_in(wire_d27_47),.data_out(wire_d27_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802749(.data_in(wire_d27_48),.data_out(wire_d27_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802750(.data_in(wire_d27_49),.data_out(wire_d27_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802751(.data_in(wire_d27_50),.data_out(wire_d27_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802752(.data_in(wire_d27_51),.data_out(wire_d27_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802753(.data_in(wire_d27_52),.data_out(wire_d27_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802754(.data_in(wire_d27_53),.data_out(wire_d27_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802755(.data_in(wire_d27_54),.data_out(wire_d27_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802756(.data_in(wire_d27_55),.data_out(wire_d27_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802757(.data_in(wire_d27_56),.data_out(wire_d27_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802758(.data_in(wire_d27_57),.data_out(wire_d27_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802759(.data_in(wire_d27_58),.data_out(wire_d27_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802760(.data_in(wire_d27_59),.data_out(wire_d27_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802761(.data_in(wire_d27_60),.data_out(wire_d27_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802762(.data_in(wire_d27_61),.data_out(wire_d27_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802763(.data_in(wire_d27_62),.data_out(wire_d27_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802764(.data_in(wire_d27_63),.data_out(wire_d27_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802765(.data_in(wire_d27_64),.data_out(wire_d27_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802766(.data_in(wire_d27_65),.data_out(wire_d27_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802767(.data_in(wire_d27_66),.data_out(wire_d27_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802768(.data_in(wire_d27_67),.data_out(wire_d27_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802769(.data_in(wire_d27_68),.data_out(wire_d27_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802770(.data_in(wire_d27_69),.data_out(wire_d27_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802771(.data_in(wire_d27_70),.data_out(wire_d27_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802772(.data_in(wire_d27_71),.data_out(wire_d27_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802773(.data_in(wire_d27_72),.data_out(wire_d27_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802774(.data_in(wire_d27_73),.data_out(wire_d27_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802775(.data_in(wire_d27_74),.data_out(wire_d27_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802776(.data_in(wire_d27_75),.data_out(wire_d27_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802777(.data_in(wire_d27_76),.data_out(wire_d27_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802778(.data_in(wire_d27_77),.data_out(wire_d27_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802779(.data_in(wire_d27_78),.data_out(d_out27),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance290280(.data_in(d_in28),.data_out(wire_d28_0),.clk(clk),.rst(rst));            //channel 29
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance290281(.data_in(wire_d28_0),.data_out(wire_d28_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance290282(.data_in(wire_d28_1),.data_out(wire_d28_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance290283(.data_in(wire_d28_2),.data_out(wire_d28_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance290284(.data_in(wire_d28_3),.data_out(wire_d28_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance290285(.data_in(wire_d28_4),.data_out(wire_d28_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance290286(.data_in(wire_d28_5),.data_out(wire_d28_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance290287(.data_in(wire_d28_6),.data_out(wire_d28_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance290288(.data_in(wire_d28_7),.data_out(wire_d28_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance290289(.data_in(wire_d28_8),.data_out(wire_d28_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902810(.data_in(wire_d28_9),.data_out(wire_d28_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902811(.data_in(wire_d28_10),.data_out(wire_d28_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902812(.data_in(wire_d28_11),.data_out(wire_d28_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902813(.data_in(wire_d28_12),.data_out(wire_d28_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902814(.data_in(wire_d28_13),.data_out(wire_d28_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902815(.data_in(wire_d28_14),.data_out(wire_d28_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902816(.data_in(wire_d28_15),.data_out(wire_d28_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902817(.data_in(wire_d28_16),.data_out(wire_d28_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902818(.data_in(wire_d28_17),.data_out(wire_d28_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902819(.data_in(wire_d28_18),.data_out(wire_d28_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902820(.data_in(wire_d28_19),.data_out(wire_d28_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902821(.data_in(wire_d28_20),.data_out(wire_d28_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902822(.data_in(wire_d28_21),.data_out(wire_d28_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902823(.data_in(wire_d28_22),.data_out(wire_d28_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902824(.data_in(wire_d28_23),.data_out(wire_d28_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902825(.data_in(wire_d28_24),.data_out(wire_d28_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902826(.data_in(wire_d28_25),.data_out(wire_d28_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902827(.data_in(wire_d28_26),.data_out(wire_d28_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902828(.data_in(wire_d28_27),.data_out(wire_d28_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902829(.data_in(wire_d28_28),.data_out(wire_d28_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902830(.data_in(wire_d28_29),.data_out(wire_d28_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902831(.data_in(wire_d28_30),.data_out(wire_d28_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902832(.data_in(wire_d28_31),.data_out(wire_d28_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902833(.data_in(wire_d28_32),.data_out(wire_d28_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902834(.data_in(wire_d28_33),.data_out(wire_d28_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902835(.data_in(wire_d28_34),.data_out(wire_d28_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902836(.data_in(wire_d28_35),.data_out(wire_d28_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902837(.data_in(wire_d28_36),.data_out(wire_d28_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902838(.data_in(wire_d28_37),.data_out(wire_d28_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902839(.data_in(wire_d28_38),.data_out(wire_d28_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902840(.data_in(wire_d28_39),.data_out(wire_d28_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902841(.data_in(wire_d28_40),.data_out(wire_d28_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902842(.data_in(wire_d28_41),.data_out(wire_d28_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902843(.data_in(wire_d28_42),.data_out(wire_d28_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902844(.data_in(wire_d28_43),.data_out(wire_d28_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902845(.data_in(wire_d28_44),.data_out(wire_d28_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902846(.data_in(wire_d28_45),.data_out(wire_d28_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902847(.data_in(wire_d28_46),.data_out(wire_d28_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902848(.data_in(wire_d28_47),.data_out(wire_d28_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902849(.data_in(wire_d28_48),.data_out(wire_d28_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902850(.data_in(wire_d28_49),.data_out(wire_d28_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902851(.data_in(wire_d28_50),.data_out(wire_d28_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902852(.data_in(wire_d28_51),.data_out(wire_d28_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902853(.data_in(wire_d28_52),.data_out(wire_d28_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902854(.data_in(wire_d28_53),.data_out(wire_d28_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902855(.data_in(wire_d28_54),.data_out(wire_d28_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902856(.data_in(wire_d28_55),.data_out(wire_d28_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902857(.data_in(wire_d28_56),.data_out(wire_d28_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902858(.data_in(wire_d28_57),.data_out(wire_d28_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902859(.data_in(wire_d28_58),.data_out(wire_d28_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902860(.data_in(wire_d28_59),.data_out(wire_d28_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902861(.data_in(wire_d28_60),.data_out(wire_d28_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902862(.data_in(wire_d28_61),.data_out(wire_d28_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902863(.data_in(wire_d28_62),.data_out(wire_d28_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902864(.data_in(wire_d28_63),.data_out(wire_d28_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902865(.data_in(wire_d28_64),.data_out(wire_d28_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902866(.data_in(wire_d28_65),.data_out(wire_d28_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902867(.data_in(wire_d28_66),.data_out(wire_d28_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902868(.data_in(wire_d28_67),.data_out(wire_d28_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902869(.data_in(wire_d28_68),.data_out(wire_d28_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902870(.data_in(wire_d28_69),.data_out(wire_d28_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902871(.data_in(wire_d28_70),.data_out(wire_d28_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902872(.data_in(wire_d28_71),.data_out(wire_d28_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902873(.data_in(wire_d28_72),.data_out(wire_d28_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902874(.data_in(wire_d28_73),.data_out(wire_d28_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902875(.data_in(wire_d28_74),.data_out(wire_d28_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902876(.data_in(wire_d28_75),.data_out(wire_d28_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902877(.data_in(wire_d28_76),.data_out(wire_d28_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902878(.data_in(wire_d28_77),.data_out(wire_d28_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902879(.data_in(wire_d28_78),.data_out(d_out28),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance300290(.data_in(d_in29),.data_out(wire_d29_0),.clk(clk),.rst(rst));            //channel 30
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance300291(.data_in(wire_d29_0),.data_out(wire_d29_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance300292(.data_in(wire_d29_1),.data_out(wire_d29_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance300293(.data_in(wire_d29_2),.data_out(wire_d29_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance300294(.data_in(wire_d29_3),.data_out(wire_d29_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance300295(.data_in(wire_d29_4),.data_out(wire_d29_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance300296(.data_in(wire_d29_5),.data_out(wire_d29_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance300297(.data_in(wire_d29_6),.data_out(wire_d29_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance300298(.data_in(wire_d29_7),.data_out(wire_d29_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance300299(.data_in(wire_d29_8),.data_out(wire_d29_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002910(.data_in(wire_d29_9),.data_out(wire_d29_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002911(.data_in(wire_d29_10),.data_out(wire_d29_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002912(.data_in(wire_d29_11),.data_out(wire_d29_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002913(.data_in(wire_d29_12),.data_out(wire_d29_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002914(.data_in(wire_d29_13),.data_out(wire_d29_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002915(.data_in(wire_d29_14),.data_out(wire_d29_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002916(.data_in(wire_d29_15),.data_out(wire_d29_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002917(.data_in(wire_d29_16),.data_out(wire_d29_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002918(.data_in(wire_d29_17),.data_out(wire_d29_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002919(.data_in(wire_d29_18),.data_out(wire_d29_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002920(.data_in(wire_d29_19),.data_out(wire_d29_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002921(.data_in(wire_d29_20),.data_out(wire_d29_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002922(.data_in(wire_d29_21),.data_out(wire_d29_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002923(.data_in(wire_d29_22),.data_out(wire_d29_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002924(.data_in(wire_d29_23),.data_out(wire_d29_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002925(.data_in(wire_d29_24),.data_out(wire_d29_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002926(.data_in(wire_d29_25),.data_out(wire_d29_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002927(.data_in(wire_d29_26),.data_out(wire_d29_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002928(.data_in(wire_d29_27),.data_out(wire_d29_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002929(.data_in(wire_d29_28),.data_out(wire_d29_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002930(.data_in(wire_d29_29),.data_out(wire_d29_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002931(.data_in(wire_d29_30),.data_out(wire_d29_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002932(.data_in(wire_d29_31),.data_out(wire_d29_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002933(.data_in(wire_d29_32),.data_out(wire_d29_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002934(.data_in(wire_d29_33),.data_out(wire_d29_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002935(.data_in(wire_d29_34),.data_out(wire_d29_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002936(.data_in(wire_d29_35),.data_out(wire_d29_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002937(.data_in(wire_d29_36),.data_out(wire_d29_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002938(.data_in(wire_d29_37),.data_out(wire_d29_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002939(.data_in(wire_d29_38),.data_out(wire_d29_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002940(.data_in(wire_d29_39),.data_out(wire_d29_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002941(.data_in(wire_d29_40),.data_out(wire_d29_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002942(.data_in(wire_d29_41),.data_out(wire_d29_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002943(.data_in(wire_d29_42),.data_out(wire_d29_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002944(.data_in(wire_d29_43),.data_out(wire_d29_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002945(.data_in(wire_d29_44),.data_out(wire_d29_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002946(.data_in(wire_d29_45),.data_out(wire_d29_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002947(.data_in(wire_d29_46),.data_out(wire_d29_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002948(.data_in(wire_d29_47),.data_out(wire_d29_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002949(.data_in(wire_d29_48),.data_out(wire_d29_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002950(.data_in(wire_d29_49),.data_out(wire_d29_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002951(.data_in(wire_d29_50),.data_out(wire_d29_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002952(.data_in(wire_d29_51),.data_out(wire_d29_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002953(.data_in(wire_d29_52),.data_out(wire_d29_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002954(.data_in(wire_d29_53),.data_out(wire_d29_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002955(.data_in(wire_d29_54),.data_out(wire_d29_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002956(.data_in(wire_d29_55),.data_out(wire_d29_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002957(.data_in(wire_d29_56),.data_out(wire_d29_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002958(.data_in(wire_d29_57),.data_out(wire_d29_58),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002959(.data_in(wire_d29_58),.data_out(wire_d29_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002960(.data_in(wire_d29_59),.data_out(wire_d29_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002961(.data_in(wire_d29_60),.data_out(wire_d29_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002962(.data_in(wire_d29_61),.data_out(wire_d29_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002963(.data_in(wire_d29_62),.data_out(wire_d29_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002964(.data_in(wire_d29_63),.data_out(wire_d29_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002965(.data_in(wire_d29_64),.data_out(wire_d29_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002966(.data_in(wire_d29_65),.data_out(wire_d29_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002967(.data_in(wire_d29_66),.data_out(wire_d29_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002968(.data_in(wire_d29_67),.data_out(wire_d29_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002969(.data_in(wire_d29_68),.data_out(wire_d29_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002970(.data_in(wire_d29_69),.data_out(wire_d29_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002971(.data_in(wire_d29_70),.data_out(wire_d29_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002972(.data_in(wire_d29_71),.data_out(wire_d29_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002973(.data_in(wire_d29_72),.data_out(wire_d29_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002974(.data_in(wire_d29_73),.data_out(wire_d29_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002975(.data_in(wire_d29_74),.data_out(wire_d29_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002976(.data_in(wire_d29_75),.data_out(wire_d29_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002977(.data_in(wire_d29_76),.data_out(wire_d29_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002978(.data_in(wire_d29_77),.data_out(wire_d29_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002979(.data_in(wire_d29_78),.data_out(d_out29),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance310300(.data_in(d_in30),.data_out(wire_d30_0),.clk(clk),.rst(rst));            //channel 31
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance310301(.data_in(wire_d30_0),.data_out(wire_d30_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance310302(.data_in(wire_d30_1),.data_out(wire_d30_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance310303(.data_in(wire_d30_2),.data_out(wire_d30_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance310304(.data_in(wire_d30_3),.data_out(wire_d30_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance310305(.data_in(wire_d30_4),.data_out(wire_d30_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance310306(.data_in(wire_d30_5),.data_out(wire_d30_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance310307(.data_in(wire_d30_6),.data_out(wire_d30_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance310308(.data_in(wire_d30_7),.data_out(wire_d30_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance310309(.data_in(wire_d30_8),.data_out(wire_d30_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103010(.data_in(wire_d30_9),.data_out(wire_d30_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103011(.data_in(wire_d30_10),.data_out(wire_d30_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103012(.data_in(wire_d30_11),.data_out(wire_d30_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103013(.data_in(wire_d30_12),.data_out(wire_d30_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103014(.data_in(wire_d30_13),.data_out(wire_d30_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103015(.data_in(wire_d30_14),.data_out(wire_d30_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103016(.data_in(wire_d30_15),.data_out(wire_d30_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103017(.data_in(wire_d30_16),.data_out(wire_d30_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103018(.data_in(wire_d30_17),.data_out(wire_d30_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103019(.data_in(wire_d30_18),.data_out(wire_d30_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103020(.data_in(wire_d30_19),.data_out(wire_d30_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103021(.data_in(wire_d30_20),.data_out(wire_d30_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103022(.data_in(wire_d30_21),.data_out(wire_d30_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103023(.data_in(wire_d30_22),.data_out(wire_d30_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103024(.data_in(wire_d30_23),.data_out(wire_d30_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103025(.data_in(wire_d30_24),.data_out(wire_d30_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103026(.data_in(wire_d30_25),.data_out(wire_d30_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103027(.data_in(wire_d30_26),.data_out(wire_d30_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103028(.data_in(wire_d30_27),.data_out(wire_d30_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103029(.data_in(wire_d30_28),.data_out(wire_d30_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103030(.data_in(wire_d30_29),.data_out(wire_d30_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103031(.data_in(wire_d30_30),.data_out(wire_d30_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103032(.data_in(wire_d30_31),.data_out(wire_d30_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103033(.data_in(wire_d30_32),.data_out(wire_d30_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103034(.data_in(wire_d30_33),.data_out(wire_d30_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103035(.data_in(wire_d30_34),.data_out(wire_d30_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103036(.data_in(wire_d30_35),.data_out(wire_d30_36),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103037(.data_in(wire_d30_36),.data_out(wire_d30_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103038(.data_in(wire_d30_37),.data_out(wire_d30_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103039(.data_in(wire_d30_38),.data_out(wire_d30_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103040(.data_in(wire_d30_39),.data_out(wire_d30_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103041(.data_in(wire_d30_40),.data_out(wire_d30_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103042(.data_in(wire_d30_41),.data_out(wire_d30_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103043(.data_in(wire_d30_42),.data_out(wire_d30_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103044(.data_in(wire_d30_43),.data_out(wire_d30_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103045(.data_in(wire_d30_44),.data_out(wire_d30_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103046(.data_in(wire_d30_45),.data_out(wire_d30_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103047(.data_in(wire_d30_46),.data_out(wire_d30_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103048(.data_in(wire_d30_47),.data_out(wire_d30_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103049(.data_in(wire_d30_48),.data_out(wire_d30_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103050(.data_in(wire_d30_49),.data_out(wire_d30_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103051(.data_in(wire_d30_50),.data_out(wire_d30_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103052(.data_in(wire_d30_51),.data_out(wire_d30_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103053(.data_in(wire_d30_52),.data_out(wire_d30_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103054(.data_in(wire_d30_53),.data_out(wire_d30_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103055(.data_in(wire_d30_54),.data_out(wire_d30_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103056(.data_in(wire_d30_55),.data_out(wire_d30_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103057(.data_in(wire_d30_56),.data_out(wire_d30_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103058(.data_in(wire_d30_57),.data_out(wire_d30_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103059(.data_in(wire_d30_58),.data_out(wire_d30_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103060(.data_in(wire_d30_59),.data_out(wire_d30_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103061(.data_in(wire_d30_60),.data_out(wire_d30_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103062(.data_in(wire_d30_61),.data_out(wire_d30_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103063(.data_in(wire_d30_62),.data_out(wire_d30_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103064(.data_in(wire_d30_63),.data_out(wire_d30_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103065(.data_in(wire_d30_64),.data_out(wire_d30_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103066(.data_in(wire_d30_65),.data_out(wire_d30_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103067(.data_in(wire_d30_66),.data_out(wire_d30_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103068(.data_in(wire_d30_67),.data_out(wire_d30_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103069(.data_in(wire_d30_68),.data_out(wire_d30_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103070(.data_in(wire_d30_69),.data_out(wire_d30_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103071(.data_in(wire_d30_70),.data_out(wire_d30_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103072(.data_in(wire_d30_71),.data_out(wire_d30_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103073(.data_in(wire_d30_72),.data_out(wire_d30_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103074(.data_in(wire_d30_73),.data_out(wire_d30_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103075(.data_in(wire_d30_74),.data_out(wire_d30_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103076(.data_in(wire_d30_75),.data_out(wire_d30_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103077(.data_in(wire_d30_76),.data_out(wire_d30_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103078(.data_in(wire_d30_77),.data_out(wire_d30_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103079(.data_in(wire_d30_78),.data_out(d_out30),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance320310(.data_in(d_in31),.data_out(wire_d31_0),.clk(clk),.rst(rst));            //channel 32
	encoder #(.WIDTH(WIDTH)) encoder_instance320311(.data_in(wire_d31_0),.data_out(wire_d31_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance320312(.data_in(wire_d31_1),.data_out(wire_d31_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance320313(.data_in(wire_d31_2),.data_out(wire_d31_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance320314(.data_in(wire_d31_3),.data_out(wire_d31_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance320315(.data_in(wire_d31_4),.data_out(wire_d31_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance320316(.data_in(wire_d31_5),.data_out(wire_d31_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance320317(.data_in(wire_d31_6),.data_out(wire_d31_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance320318(.data_in(wire_d31_7),.data_out(wire_d31_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance320319(.data_in(wire_d31_8),.data_out(wire_d31_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203110(.data_in(wire_d31_9),.data_out(wire_d31_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203111(.data_in(wire_d31_10),.data_out(wire_d31_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203112(.data_in(wire_d31_11),.data_out(wire_d31_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203113(.data_in(wire_d31_12),.data_out(wire_d31_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203114(.data_in(wire_d31_13),.data_out(wire_d31_14),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203115(.data_in(wire_d31_14),.data_out(wire_d31_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203116(.data_in(wire_d31_15),.data_out(wire_d31_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203117(.data_in(wire_d31_16),.data_out(wire_d31_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203118(.data_in(wire_d31_17),.data_out(wire_d31_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203119(.data_in(wire_d31_18),.data_out(wire_d31_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203120(.data_in(wire_d31_19),.data_out(wire_d31_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203121(.data_in(wire_d31_20),.data_out(wire_d31_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203122(.data_in(wire_d31_21),.data_out(wire_d31_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203123(.data_in(wire_d31_22),.data_out(wire_d31_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203124(.data_in(wire_d31_23),.data_out(wire_d31_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203125(.data_in(wire_d31_24),.data_out(wire_d31_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203126(.data_in(wire_d31_25),.data_out(wire_d31_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203127(.data_in(wire_d31_26),.data_out(wire_d31_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203128(.data_in(wire_d31_27),.data_out(wire_d31_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203129(.data_in(wire_d31_28),.data_out(wire_d31_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203130(.data_in(wire_d31_29),.data_out(wire_d31_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203131(.data_in(wire_d31_30),.data_out(wire_d31_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203132(.data_in(wire_d31_31),.data_out(wire_d31_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203133(.data_in(wire_d31_32),.data_out(wire_d31_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203134(.data_in(wire_d31_33),.data_out(wire_d31_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203135(.data_in(wire_d31_34),.data_out(wire_d31_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203136(.data_in(wire_d31_35),.data_out(wire_d31_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203137(.data_in(wire_d31_36),.data_out(wire_d31_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203138(.data_in(wire_d31_37),.data_out(wire_d31_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203139(.data_in(wire_d31_38),.data_out(wire_d31_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203140(.data_in(wire_d31_39),.data_out(wire_d31_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203141(.data_in(wire_d31_40),.data_out(wire_d31_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203142(.data_in(wire_d31_41),.data_out(wire_d31_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203143(.data_in(wire_d31_42),.data_out(wire_d31_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203144(.data_in(wire_d31_43),.data_out(wire_d31_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203145(.data_in(wire_d31_44),.data_out(wire_d31_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203146(.data_in(wire_d31_45),.data_out(wire_d31_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203147(.data_in(wire_d31_46),.data_out(wire_d31_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203148(.data_in(wire_d31_47),.data_out(wire_d31_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203149(.data_in(wire_d31_48),.data_out(wire_d31_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203150(.data_in(wire_d31_49),.data_out(wire_d31_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203151(.data_in(wire_d31_50),.data_out(wire_d31_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203152(.data_in(wire_d31_51),.data_out(wire_d31_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203153(.data_in(wire_d31_52),.data_out(wire_d31_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203154(.data_in(wire_d31_53),.data_out(wire_d31_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203155(.data_in(wire_d31_54),.data_out(wire_d31_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203156(.data_in(wire_d31_55),.data_out(wire_d31_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203157(.data_in(wire_d31_56),.data_out(wire_d31_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203158(.data_in(wire_d31_57),.data_out(wire_d31_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203159(.data_in(wire_d31_58),.data_out(wire_d31_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203160(.data_in(wire_d31_59),.data_out(wire_d31_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203161(.data_in(wire_d31_60),.data_out(wire_d31_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203162(.data_in(wire_d31_61),.data_out(wire_d31_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203163(.data_in(wire_d31_62),.data_out(wire_d31_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203164(.data_in(wire_d31_63),.data_out(wire_d31_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203165(.data_in(wire_d31_64),.data_out(wire_d31_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203166(.data_in(wire_d31_65),.data_out(wire_d31_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203167(.data_in(wire_d31_66),.data_out(wire_d31_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203168(.data_in(wire_d31_67),.data_out(wire_d31_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203169(.data_in(wire_d31_68),.data_out(wire_d31_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203170(.data_in(wire_d31_69),.data_out(wire_d31_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203171(.data_in(wire_d31_70),.data_out(wire_d31_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203172(.data_in(wire_d31_71),.data_out(wire_d31_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203173(.data_in(wire_d31_72),.data_out(wire_d31_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203174(.data_in(wire_d31_73),.data_out(wire_d31_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203175(.data_in(wire_d31_74),.data_out(wire_d31_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203176(.data_in(wire_d31_75),.data_out(wire_d31_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203177(.data_in(wire_d31_76),.data_out(wire_d31_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203178(.data_in(wire_d31_77),.data_out(wire_d31_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203179(.data_in(wire_d31_78),.data_out(d_out31),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance330320(.data_in(d_in32),.data_out(wire_d32_0),.clk(clk),.rst(rst));            //channel 33
	decoder_top #(.WIDTH(WIDTH)) decoder_instance330321(.data_in(wire_d32_0),.data_out(wire_d32_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance330322(.data_in(wire_d32_1),.data_out(wire_d32_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance330323(.data_in(wire_d32_2),.data_out(wire_d32_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance330324(.data_in(wire_d32_3),.data_out(wire_d32_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance330325(.data_in(wire_d32_4),.data_out(wire_d32_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance330326(.data_in(wire_d32_5),.data_out(wire_d32_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance330327(.data_in(wire_d32_6),.data_out(wire_d32_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance330328(.data_in(wire_d32_7),.data_out(wire_d32_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance330329(.data_in(wire_d32_8),.data_out(wire_d32_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303210(.data_in(wire_d32_9),.data_out(wire_d32_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303211(.data_in(wire_d32_10),.data_out(wire_d32_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303212(.data_in(wire_d32_11),.data_out(wire_d32_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303213(.data_in(wire_d32_12),.data_out(wire_d32_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303214(.data_in(wire_d32_13),.data_out(wire_d32_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303215(.data_in(wire_d32_14),.data_out(wire_d32_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303216(.data_in(wire_d32_15),.data_out(wire_d32_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303217(.data_in(wire_d32_16),.data_out(wire_d32_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303218(.data_in(wire_d32_17),.data_out(wire_d32_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303219(.data_in(wire_d32_18),.data_out(wire_d32_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303220(.data_in(wire_d32_19),.data_out(wire_d32_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303221(.data_in(wire_d32_20),.data_out(wire_d32_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303222(.data_in(wire_d32_21),.data_out(wire_d32_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303223(.data_in(wire_d32_22),.data_out(wire_d32_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303224(.data_in(wire_d32_23),.data_out(wire_d32_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303225(.data_in(wire_d32_24),.data_out(wire_d32_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303226(.data_in(wire_d32_25),.data_out(wire_d32_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303227(.data_in(wire_d32_26),.data_out(wire_d32_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303228(.data_in(wire_d32_27),.data_out(wire_d32_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303229(.data_in(wire_d32_28),.data_out(wire_d32_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303230(.data_in(wire_d32_29),.data_out(wire_d32_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303231(.data_in(wire_d32_30),.data_out(wire_d32_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303232(.data_in(wire_d32_31),.data_out(wire_d32_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303233(.data_in(wire_d32_32),.data_out(wire_d32_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303234(.data_in(wire_d32_33),.data_out(wire_d32_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303235(.data_in(wire_d32_34),.data_out(wire_d32_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303236(.data_in(wire_d32_35),.data_out(wire_d32_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303237(.data_in(wire_d32_36),.data_out(wire_d32_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303238(.data_in(wire_d32_37),.data_out(wire_d32_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303239(.data_in(wire_d32_38),.data_out(wire_d32_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303240(.data_in(wire_d32_39),.data_out(wire_d32_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303241(.data_in(wire_d32_40),.data_out(wire_d32_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303242(.data_in(wire_d32_41),.data_out(wire_d32_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303243(.data_in(wire_d32_42),.data_out(wire_d32_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303244(.data_in(wire_d32_43),.data_out(wire_d32_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303245(.data_in(wire_d32_44),.data_out(wire_d32_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303246(.data_in(wire_d32_45),.data_out(wire_d32_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303247(.data_in(wire_d32_46),.data_out(wire_d32_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303248(.data_in(wire_d32_47),.data_out(wire_d32_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303249(.data_in(wire_d32_48),.data_out(wire_d32_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303250(.data_in(wire_d32_49),.data_out(wire_d32_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303251(.data_in(wire_d32_50),.data_out(wire_d32_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303252(.data_in(wire_d32_51),.data_out(wire_d32_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303253(.data_in(wire_d32_52),.data_out(wire_d32_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303254(.data_in(wire_d32_53),.data_out(wire_d32_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303255(.data_in(wire_d32_54),.data_out(wire_d32_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303256(.data_in(wire_d32_55),.data_out(wire_d32_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303257(.data_in(wire_d32_56),.data_out(wire_d32_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303258(.data_in(wire_d32_57),.data_out(wire_d32_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303259(.data_in(wire_d32_58),.data_out(wire_d32_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303260(.data_in(wire_d32_59),.data_out(wire_d32_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303261(.data_in(wire_d32_60),.data_out(wire_d32_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303262(.data_in(wire_d32_61),.data_out(wire_d32_62),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303263(.data_in(wire_d32_62),.data_out(wire_d32_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303264(.data_in(wire_d32_63),.data_out(wire_d32_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303265(.data_in(wire_d32_64),.data_out(wire_d32_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303266(.data_in(wire_d32_65),.data_out(wire_d32_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303267(.data_in(wire_d32_66),.data_out(wire_d32_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303268(.data_in(wire_d32_67),.data_out(wire_d32_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303269(.data_in(wire_d32_68),.data_out(wire_d32_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303270(.data_in(wire_d32_69),.data_out(wire_d32_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303271(.data_in(wire_d32_70),.data_out(wire_d32_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303272(.data_in(wire_d32_71),.data_out(wire_d32_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303273(.data_in(wire_d32_72),.data_out(wire_d32_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303274(.data_in(wire_d32_73),.data_out(wire_d32_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303275(.data_in(wire_d32_74),.data_out(wire_d32_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303276(.data_in(wire_d32_75),.data_out(wire_d32_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303277(.data_in(wire_d32_76),.data_out(wire_d32_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303278(.data_in(wire_d32_77),.data_out(wire_d32_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303279(.data_in(wire_d32_78),.data_out(d_out32),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance340330(.data_in(d_in33),.data_out(wire_d33_0),.clk(clk),.rst(rst));            //channel 34
	decoder_top #(.WIDTH(WIDTH)) decoder_instance340331(.data_in(wire_d33_0),.data_out(wire_d33_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance340332(.data_in(wire_d33_1),.data_out(wire_d33_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance340333(.data_in(wire_d33_2),.data_out(wire_d33_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance340334(.data_in(wire_d33_3),.data_out(wire_d33_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance340335(.data_in(wire_d33_4),.data_out(wire_d33_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance340336(.data_in(wire_d33_5),.data_out(wire_d33_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance340337(.data_in(wire_d33_6),.data_out(wire_d33_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance340338(.data_in(wire_d33_7),.data_out(wire_d33_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance340339(.data_in(wire_d33_8),.data_out(wire_d33_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403310(.data_in(wire_d33_9),.data_out(wire_d33_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403311(.data_in(wire_d33_10),.data_out(wire_d33_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403312(.data_in(wire_d33_11),.data_out(wire_d33_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403313(.data_in(wire_d33_12),.data_out(wire_d33_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403314(.data_in(wire_d33_13),.data_out(wire_d33_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403315(.data_in(wire_d33_14),.data_out(wire_d33_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403316(.data_in(wire_d33_15),.data_out(wire_d33_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403317(.data_in(wire_d33_16),.data_out(wire_d33_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403318(.data_in(wire_d33_17),.data_out(wire_d33_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403319(.data_in(wire_d33_18),.data_out(wire_d33_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403320(.data_in(wire_d33_19),.data_out(wire_d33_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403321(.data_in(wire_d33_20),.data_out(wire_d33_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403322(.data_in(wire_d33_21),.data_out(wire_d33_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403323(.data_in(wire_d33_22),.data_out(wire_d33_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403324(.data_in(wire_d33_23),.data_out(wire_d33_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403325(.data_in(wire_d33_24),.data_out(wire_d33_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403326(.data_in(wire_d33_25),.data_out(wire_d33_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403327(.data_in(wire_d33_26),.data_out(wire_d33_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403328(.data_in(wire_d33_27),.data_out(wire_d33_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403329(.data_in(wire_d33_28),.data_out(wire_d33_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403330(.data_in(wire_d33_29),.data_out(wire_d33_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403331(.data_in(wire_d33_30),.data_out(wire_d33_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403332(.data_in(wire_d33_31),.data_out(wire_d33_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403333(.data_in(wire_d33_32),.data_out(wire_d33_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403334(.data_in(wire_d33_33),.data_out(wire_d33_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403335(.data_in(wire_d33_34),.data_out(wire_d33_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403336(.data_in(wire_d33_35),.data_out(wire_d33_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403337(.data_in(wire_d33_36),.data_out(wire_d33_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403338(.data_in(wire_d33_37),.data_out(wire_d33_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403339(.data_in(wire_d33_38),.data_out(wire_d33_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403340(.data_in(wire_d33_39),.data_out(wire_d33_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403341(.data_in(wire_d33_40),.data_out(wire_d33_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403342(.data_in(wire_d33_41),.data_out(wire_d33_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403343(.data_in(wire_d33_42),.data_out(wire_d33_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403344(.data_in(wire_d33_43),.data_out(wire_d33_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403345(.data_in(wire_d33_44),.data_out(wire_d33_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403346(.data_in(wire_d33_45),.data_out(wire_d33_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403347(.data_in(wire_d33_46),.data_out(wire_d33_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403348(.data_in(wire_d33_47),.data_out(wire_d33_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403349(.data_in(wire_d33_48),.data_out(wire_d33_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403350(.data_in(wire_d33_49),.data_out(wire_d33_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403351(.data_in(wire_d33_50),.data_out(wire_d33_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403352(.data_in(wire_d33_51),.data_out(wire_d33_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403353(.data_in(wire_d33_52),.data_out(wire_d33_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403354(.data_in(wire_d33_53),.data_out(wire_d33_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403355(.data_in(wire_d33_54),.data_out(wire_d33_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403356(.data_in(wire_d33_55),.data_out(wire_d33_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403357(.data_in(wire_d33_56),.data_out(wire_d33_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403358(.data_in(wire_d33_57),.data_out(wire_d33_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403359(.data_in(wire_d33_58),.data_out(wire_d33_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403360(.data_in(wire_d33_59),.data_out(wire_d33_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403361(.data_in(wire_d33_60),.data_out(wire_d33_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403362(.data_in(wire_d33_61),.data_out(wire_d33_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403363(.data_in(wire_d33_62),.data_out(wire_d33_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403364(.data_in(wire_d33_63),.data_out(wire_d33_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403365(.data_in(wire_d33_64),.data_out(wire_d33_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403366(.data_in(wire_d33_65),.data_out(wire_d33_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403367(.data_in(wire_d33_66),.data_out(wire_d33_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403368(.data_in(wire_d33_67),.data_out(wire_d33_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403369(.data_in(wire_d33_68),.data_out(wire_d33_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403370(.data_in(wire_d33_69),.data_out(wire_d33_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403371(.data_in(wire_d33_70),.data_out(wire_d33_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403372(.data_in(wire_d33_71),.data_out(wire_d33_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403373(.data_in(wire_d33_72),.data_out(wire_d33_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403374(.data_in(wire_d33_73),.data_out(wire_d33_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403375(.data_in(wire_d33_74),.data_out(wire_d33_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403376(.data_in(wire_d33_75),.data_out(wire_d33_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403377(.data_in(wire_d33_76),.data_out(wire_d33_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403378(.data_in(wire_d33_77),.data_out(wire_d33_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403379(.data_in(wire_d33_78),.data_out(d_out33),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance350340(.data_in(d_in34),.data_out(wire_d34_0),.clk(clk),.rst(rst));            //channel 35
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance350341(.data_in(wire_d34_0),.data_out(wire_d34_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance350342(.data_in(wire_d34_1),.data_out(wire_d34_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance350343(.data_in(wire_d34_2),.data_out(wire_d34_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance350344(.data_in(wire_d34_3),.data_out(wire_d34_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance350345(.data_in(wire_d34_4),.data_out(wire_d34_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance350346(.data_in(wire_d34_5),.data_out(wire_d34_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance350347(.data_in(wire_d34_6),.data_out(wire_d34_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance350348(.data_in(wire_d34_7),.data_out(wire_d34_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance350349(.data_in(wire_d34_8),.data_out(wire_d34_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503410(.data_in(wire_d34_9),.data_out(wire_d34_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503411(.data_in(wire_d34_10),.data_out(wire_d34_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503412(.data_in(wire_d34_11),.data_out(wire_d34_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503413(.data_in(wire_d34_12),.data_out(wire_d34_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503414(.data_in(wire_d34_13),.data_out(wire_d34_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503415(.data_in(wire_d34_14),.data_out(wire_d34_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503416(.data_in(wire_d34_15),.data_out(wire_d34_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503417(.data_in(wire_d34_16),.data_out(wire_d34_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503418(.data_in(wire_d34_17),.data_out(wire_d34_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503419(.data_in(wire_d34_18),.data_out(wire_d34_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503420(.data_in(wire_d34_19),.data_out(wire_d34_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503421(.data_in(wire_d34_20),.data_out(wire_d34_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503422(.data_in(wire_d34_21),.data_out(wire_d34_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503423(.data_in(wire_d34_22),.data_out(wire_d34_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503424(.data_in(wire_d34_23),.data_out(wire_d34_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503425(.data_in(wire_d34_24),.data_out(wire_d34_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503426(.data_in(wire_d34_25),.data_out(wire_d34_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503427(.data_in(wire_d34_26),.data_out(wire_d34_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503428(.data_in(wire_d34_27),.data_out(wire_d34_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503429(.data_in(wire_d34_28),.data_out(wire_d34_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503430(.data_in(wire_d34_29),.data_out(wire_d34_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503431(.data_in(wire_d34_30),.data_out(wire_d34_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503432(.data_in(wire_d34_31),.data_out(wire_d34_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503433(.data_in(wire_d34_32),.data_out(wire_d34_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503434(.data_in(wire_d34_33),.data_out(wire_d34_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503435(.data_in(wire_d34_34),.data_out(wire_d34_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503436(.data_in(wire_d34_35),.data_out(wire_d34_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503437(.data_in(wire_d34_36),.data_out(wire_d34_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503438(.data_in(wire_d34_37),.data_out(wire_d34_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503439(.data_in(wire_d34_38),.data_out(wire_d34_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503440(.data_in(wire_d34_39),.data_out(wire_d34_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503441(.data_in(wire_d34_40),.data_out(wire_d34_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503442(.data_in(wire_d34_41),.data_out(wire_d34_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503443(.data_in(wire_d34_42),.data_out(wire_d34_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503444(.data_in(wire_d34_43),.data_out(wire_d34_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503445(.data_in(wire_d34_44),.data_out(wire_d34_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503446(.data_in(wire_d34_45),.data_out(wire_d34_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503447(.data_in(wire_d34_46),.data_out(wire_d34_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503448(.data_in(wire_d34_47),.data_out(wire_d34_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503449(.data_in(wire_d34_48),.data_out(wire_d34_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503450(.data_in(wire_d34_49),.data_out(wire_d34_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503451(.data_in(wire_d34_50),.data_out(wire_d34_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503452(.data_in(wire_d34_51),.data_out(wire_d34_52),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503453(.data_in(wire_d34_52),.data_out(wire_d34_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503454(.data_in(wire_d34_53),.data_out(wire_d34_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503455(.data_in(wire_d34_54),.data_out(wire_d34_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503456(.data_in(wire_d34_55),.data_out(wire_d34_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503457(.data_in(wire_d34_56),.data_out(wire_d34_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503458(.data_in(wire_d34_57),.data_out(wire_d34_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503459(.data_in(wire_d34_58),.data_out(wire_d34_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503460(.data_in(wire_d34_59),.data_out(wire_d34_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503461(.data_in(wire_d34_60),.data_out(wire_d34_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503462(.data_in(wire_d34_61),.data_out(wire_d34_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503463(.data_in(wire_d34_62),.data_out(wire_d34_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503464(.data_in(wire_d34_63),.data_out(wire_d34_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503465(.data_in(wire_d34_64),.data_out(wire_d34_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503466(.data_in(wire_d34_65),.data_out(wire_d34_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503467(.data_in(wire_d34_66),.data_out(wire_d34_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503468(.data_in(wire_d34_67),.data_out(wire_d34_68),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503469(.data_in(wire_d34_68),.data_out(wire_d34_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503470(.data_in(wire_d34_69),.data_out(wire_d34_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503471(.data_in(wire_d34_70),.data_out(wire_d34_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503472(.data_in(wire_d34_71),.data_out(wire_d34_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503473(.data_in(wire_d34_72),.data_out(wire_d34_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503474(.data_in(wire_d34_73),.data_out(wire_d34_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503475(.data_in(wire_d34_74),.data_out(wire_d34_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503476(.data_in(wire_d34_75),.data_out(wire_d34_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503477(.data_in(wire_d34_76),.data_out(wire_d34_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503478(.data_in(wire_d34_77),.data_out(wire_d34_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503479(.data_in(wire_d34_78),.data_out(d_out34),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance360350(.data_in(d_in35),.data_out(wire_d35_0),.clk(clk),.rst(rst));            //channel 36
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance360351(.data_in(wire_d35_0),.data_out(wire_d35_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance360352(.data_in(wire_d35_1),.data_out(wire_d35_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance360353(.data_in(wire_d35_2),.data_out(wire_d35_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance360354(.data_in(wire_d35_3),.data_out(wire_d35_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance360355(.data_in(wire_d35_4),.data_out(wire_d35_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance360356(.data_in(wire_d35_5),.data_out(wire_d35_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance360357(.data_in(wire_d35_6),.data_out(wire_d35_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance360358(.data_in(wire_d35_7),.data_out(wire_d35_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance360359(.data_in(wire_d35_8),.data_out(wire_d35_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603510(.data_in(wire_d35_9),.data_out(wire_d35_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603511(.data_in(wire_d35_10),.data_out(wire_d35_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603512(.data_in(wire_d35_11),.data_out(wire_d35_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603513(.data_in(wire_d35_12),.data_out(wire_d35_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603514(.data_in(wire_d35_13),.data_out(wire_d35_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603515(.data_in(wire_d35_14),.data_out(wire_d35_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603516(.data_in(wire_d35_15),.data_out(wire_d35_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603517(.data_in(wire_d35_16),.data_out(wire_d35_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603518(.data_in(wire_d35_17),.data_out(wire_d35_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603519(.data_in(wire_d35_18),.data_out(wire_d35_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603520(.data_in(wire_d35_19),.data_out(wire_d35_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603521(.data_in(wire_d35_20),.data_out(wire_d35_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603522(.data_in(wire_d35_21),.data_out(wire_d35_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603523(.data_in(wire_d35_22),.data_out(wire_d35_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603524(.data_in(wire_d35_23),.data_out(wire_d35_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603525(.data_in(wire_d35_24),.data_out(wire_d35_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603526(.data_in(wire_d35_25),.data_out(wire_d35_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603527(.data_in(wire_d35_26),.data_out(wire_d35_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603528(.data_in(wire_d35_27),.data_out(wire_d35_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603529(.data_in(wire_d35_28),.data_out(wire_d35_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603530(.data_in(wire_d35_29),.data_out(wire_d35_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603531(.data_in(wire_d35_30),.data_out(wire_d35_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603532(.data_in(wire_d35_31),.data_out(wire_d35_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603533(.data_in(wire_d35_32),.data_out(wire_d35_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603534(.data_in(wire_d35_33),.data_out(wire_d35_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603535(.data_in(wire_d35_34),.data_out(wire_d35_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603536(.data_in(wire_d35_35),.data_out(wire_d35_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603537(.data_in(wire_d35_36),.data_out(wire_d35_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603538(.data_in(wire_d35_37),.data_out(wire_d35_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603539(.data_in(wire_d35_38),.data_out(wire_d35_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603540(.data_in(wire_d35_39),.data_out(wire_d35_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603541(.data_in(wire_d35_40),.data_out(wire_d35_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603542(.data_in(wire_d35_41),.data_out(wire_d35_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603543(.data_in(wire_d35_42),.data_out(wire_d35_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603544(.data_in(wire_d35_43),.data_out(wire_d35_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603545(.data_in(wire_d35_44),.data_out(wire_d35_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603546(.data_in(wire_d35_45),.data_out(wire_d35_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603547(.data_in(wire_d35_46),.data_out(wire_d35_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603548(.data_in(wire_d35_47),.data_out(wire_d35_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603549(.data_in(wire_d35_48),.data_out(wire_d35_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603550(.data_in(wire_d35_49),.data_out(wire_d35_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603551(.data_in(wire_d35_50),.data_out(wire_d35_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603552(.data_in(wire_d35_51),.data_out(wire_d35_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603553(.data_in(wire_d35_52),.data_out(wire_d35_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603554(.data_in(wire_d35_53),.data_out(wire_d35_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603555(.data_in(wire_d35_54),.data_out(wire_d35_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603556(.data_in(wire_d35_55),.data_out(wire_d35_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603557(.data_in(wire_d35_56),.data_out(wire_d35_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3603558(.data_in(wire_d35_57),.data_out(wire_d35_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603559(.data_in(wire_d35_58),.data_out(wire_d35_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3603560(.data_in(wire_d35_59),.data_out(wire_d35_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603561(.data_in(wire_d35_60),.data_out(wire_d35_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603562(.data_in(wire_d35_61),.data_out(wire_d35_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603563(.data_in(wire_d35_62),.data_out(wire_d35_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603564(.data_in(wire_d35_63),.data_out(wire_d35_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603565(.data_in(wire_d35_64),.data_out(wire_d35_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603566(.data_in(wire_d35_65),.data_out(wire_d35_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603567(.data_in(wire_d35_66),.data_out(wire_d35_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603568(.data_in(wire_d35_67),.data_out(wire_d35_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603569(.data_in(wire_d35_68),.data_out(wire_d35_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603570(.data_in(wire_d35_69),.data_out(wire_d35_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603571(.data_in(wire_d35_70),.data_out(wire_d35_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603572(.data_in(wire_d35_71),.data_out(wire_d35_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603573(.data_in(wire_d35_72),.data_out(wire_d35_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603574(.data_in(wire_d35_73),.data_out(wire_d35_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603575(.data_in(wire_d35_74),.data_out(wire_d35_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603576(.data_in(wire_d35_75),.data_out(wire_d35_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603577(.data_in(wire_d35_76),.data_out(wire_d35_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603578(.data_in(wire_d35_77),.data_out(wire_d35_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603579(.data_in(wire_d35_78),.data_out(d_out35),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance370360(.data_in(d_in36),.data_out(wire_d36_0),.clk(clk),.rst(rst));            //channel 37
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance370361(.data_in(wire_d36_0),.data_out(wire_d36_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance370362(.data_in(wire_d36_1),.data_out(wire_d36_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance370363(.data_in(wire_d36_2),.data_out(wire_d36_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance370364(.data_in(wire_d36_3),.data_out(wire_d36_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance370365(.data_in(wire_d36_4),.data_out(wire_d36_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance370366(.data_in(wire_d36_5),.data_out(wire_d36_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance370367(.data_in(wire_d36_6),.data_out(wire_d36_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance370368(.data_in(wire_d36_7),.data_out(wire_d36_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance370369(.data_in(wire_d36_8),.data_out(wire_d36_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703610(.data_in(wire_d36_9),.data_out(wire_d36_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703611(.data_in(wire_d36_10),.data_out(wire_d36_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703612(.data_in(wire_d36_11),.data_out(wire_d36_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703613(.data_in(wire_d36_12),.data_out(wire_d36_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703614(.data_in(wire_d36_13),.data_out(wire_d36_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703615(.data_in(wire_d36_14),.data_out(wire_d36_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703616(.data_in(wire_d36_15),.data_out(wire_d36_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703617(.data_in(wire_d36_16),.data_out(wire_d36_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703618(.data_in(wire_d36_17),.data_out(wire_d36_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703619(.data_in(wire_d36_18),.data_out(wire_d36_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703620(.data_in(wire_d36_19),.data_out(wire_d36_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703621(.data_in(wire_d36_20),.data_out(wire_d36_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703622(.data_in(wire_d36_21),.data_out(wire_d36_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703623(.data_in(wire_d36_22),.data_out(wire_d36_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703624(.data_in(wire_d36_23),.data_out(wire_d36_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703625(.data_in(wire_d36_24),.data_out(wire_d36_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703626(.data_in(wire_d36_25),.data_out(wire_d36_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703627(.data_in(wire_d36_26),.data_out(wire_d36_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703628(.data_in(wire_d36_27),.data_out(wire_d36_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703629(.data_in(wire_d36_28),.data_out(wire_d36_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703630(.data_in(wire_d36_29),.data_out(wire_d36_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703631(.data_in(wire_d36_30),.data_out(wire_d36_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703632(.data_in(wire_d36_31),.data_out(wire_d36_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703633(.data_in(wire_d36_32),.data_out(wire_d36_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703634(.data_in(wire_d36_33),.data_out(wire_d36_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703635(.data_in(wire_d36_34),.data_out(wire_d36_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703636(.data_in(wire_d36_35),.data_out(wire_d36_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703637(.data_in(wire_d36_36),.data_out(wire_d36_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703638(.data_in(wire_d36_37),.data_out(wire_d36_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703639(.data_in(wire_d36_38),.data_out(wire_d36_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703640(.data_in(wire_d36_39),.data_out(wire_d36_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703641(.data_in(wire_d36_40),.data_out(wire_d36_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703642(.data_in(wire_d36_41),.data_out(wire_d36_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703643(.data_in(wire_d36_42),.data_out(wire_d36_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703644(.data_in(wire_d36_43),.data_out(wire_d36_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703645(.data_in(wire_d36_44),.data_out(wire_d36_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703646(.data_in(wire_d36_45),.data_out(wire_d36_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703647(.data_in(wire_d36_46),.data_out(wire_d36_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703648(.data_in(wire_d36_47),.data_out(wire_d36_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703649(.data_in(wire_d36_48),.data_out(wire_d36_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703650(.data_in(wire_d36_49),.data_out(wire_d36_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703651(.data_in(wire_d36_50),.data_out(wire_d36_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703652(.data_in(wire_d36_51),.data_out(wire_d36_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703653(.data_in(wire_d36_52),.data_out(wire_d36_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703654(.data_in(wire_d36_53),.data_out(wire_d36_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703655(.data_in(wire_d36_54),.data_out(wire_d36_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703656(.data_in(wire_d36_55),.data_out(wire_d36_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703657(.data_in(wire_d36_56),.data_out(wire_d36_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703658(.data_in(wire_d36_57),.data_out(wire_d36_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703659(.data_in(wire_d36_58),.data_out(wire_d36_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703660(.data_in(wire_d36_59),.data_out(wire_d36_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703661(.data_in(wire_d36_60),.data_out(wire_d36_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703662(.data_in(wire_d36_61),.data_out(wire_d36_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703663(.data_in(wire_d36_62),.data_out(wire_d36_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703664(.data_in(wire_d36_63),.data_out(wire_d36_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703665(.data_in(wire_d36_64),.data_out(wire_d36_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703666(.data_in(wire_d36_65),.data_out(wire_d36_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703667(.data_in(wire_d36_66),.data_out(wire_d36_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703668(.data_in(wire_d36_67),.data_out(wire_d36_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703669(.data_in(wire_d36_68),.data_out(wire_d36_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703670(.data_in(wire_d36_69),.data_out(wire_d36_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703671(.data_in(wire_d36_70),.data_out(wire_d36_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703672(.data_in(wire_d36_71),.data_out(wire_d36_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703673(.data_in(wire_d36_72),.data_out(wire_d36_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703674(.data_in(wire_d36_73),.data_out(wire_d36_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703675(.data_in(wire_d36_74),.data_out(wire_d36_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703676(.data_in(wire_d36_75),.data_out(wire_d36_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703677(.data_in(wire_d36_76),.data_out(wire_d36_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703678(.data_in(wire_d36_77),.data_out(wire_d36_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703679(.data_in(wire_d36_78),.data_out(d_out36),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance380370(.data_in(d_in37),.data_out(wire_d37_0),.clk(clk),.rst(rst));            //channel 38
	invertion #(.WIDTH(WIDTH)) invertion_instance380371(.data_in(wire_d37_0),.data_out(wire_d37_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance380372(.data_in(wire_d37_1),.data_out(wire_d37_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance380373(.data_in(wire_d37_2),.data_out(wire_d37_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance380374(.data_in(wire_d37_3),.data_out(wire_d37_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance380375(.data_in(wire_d37_4),.data_out(wire_d37_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance380376(.data_in(wire_d37_5),.data_out(wire_d37_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance380377(.data_in(wire_d37_6),.data_out(wire_d37_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance380378(.data_in(wire_d37_7),.data_out(wire_d37_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance380379(.data_in(wire_d37_8),.data_out(wire_d37_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803710(.data_in(wire_d37_9),.data_out(wire_d37_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803711(.data_in(wire_d37_10),.data_out(wire_d37_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803712(.data_in(wire_d37_11),.data_out(wire_d37_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803713(.data_in(wire_d37_12),.data_out(wire_d37_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803714(.data_in(wire_d37_13),.data_out(wire_d37_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803715(.data_in(wire_d37_14),.data_out(wire_d37_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803716(.data_in(wire_d37_15),.data_out(wire_d37_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803717(.data_in(wire_d37_16),.data_out(wire_d37_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803718(.data_in(wire_d37_17),.data_out(wire_d37_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803719(.data_in(wire_d37_18),.data_out(wire_d37_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803720(.data_in(wire_d37_19),.data_out(wire_d37_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803721(.data_in(wire_d37_20),.data_out(wire_d37_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803722(.data_in(wire_d37_21),.data_out(wire_d37_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803723(.data_in(wire_d37_22),.data_out(wire_d37_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803724(.data_in(wire_d37_23),.data_out(wire_d37_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803725(.data_in(wire_d37_24),.data_out(wire_d37_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803726(.data_in(wire_d37_25),.data_out(wire_d37_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803727(.data_in(wire_d37_26),.data_out(wire_d37_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803728(.data_in(wire_d37_27),.data_out(wire_d37_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803729(.data_in(wire_d37_28),.data_out(wire_d37_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803730(.data_in(wire_d37_29),.data_out(wire_d37_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803731(.data_in(wire_d37_30),.data_out(wire_d37_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803732(.data_in(wire_d37_31),.data_out(wire_d37_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803733(.data_in(wire_d37_32),.data_out(wire_d37_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803734(.data_in(wire_d37_33),.data_out(wire_d37_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803735(.data_in(wire_d37_34),.data_out(wire_d37_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803736(.data_in(wire_d37_35),.data_out(wire_d37_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803737(.data_in(wire_d37_36),.data_out(wire_d37_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803738(.data_in(wire_d37_37),.data_out(wire_d37_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803739(.data_in(wire_d37_38),.data_out(wire_d37_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803740(.data_in(wire_d37_39),.data_out(wire_d37_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803741(.data_in(wire_d37_40),.data_out(wire_d37_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803742(.data_in(wire_d37_41),.data_out(wire_d37_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803743(.data_in(wire_d37_42),.data_out(wire_d37_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803744(.data_in(wire_d37_43),.data_out(wire_d37_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803745(.data_in(wire_d37_44),.data_out(wire_d37_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803746(.data_in(wire_d37_45),.data_out(wire_d37_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803747(.data_in(wire_d37_46),.data_out(wire_d37_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803748(.data_in(wire_d37_47),.data_out(wire_d37_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803749(.data_in(wire_d37_48),.data_out(wire_d37_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803750(.data_in(wire_d37_49),.data_out(wire_d37_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803751(.data_in(wire_d37_50),.data_out(wire_d37_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803752(.data_in(wire_d37_51),.data_out(wire_d37_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803753(.data_in(wire_d37_52),.data_out(wire_d37_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803754(.data_in(wire_d37_53),.data_out(wire_d37_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803755(.data_in(wire_d37_54),.data_out(wire_d37_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803756(.data_in(wire_d37_55),.data_out(wire_d37_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803757(.data_in(wire_d37_56),.data_out(wire_d37_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803758(.data_in(wire_d37_57),.data_out(wire_d37_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803759(.data_in(wire_d37_58),.data_out(wire_d37_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803760(.data_in(wire_d37_59),.data_out(wire_d37_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803761(.data_in(wire_d37_60),.data_out(wire_d37_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803762(.data_in(wire_d37_61),.data_out(wire_d37_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803763(.data_in(wire_d37_62),.data_out(wire_d37_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803764(.data_in(wire_d37_63),.data_out(wire_d37_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803765(.data_in(wire_d37_64),.data_out(wire_d37_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803766(.data_in(wire_d37_65),.data_out(wire_d37_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803767(.data_in(wire_d37_66),.data_out(wire_d37_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803768(.data_in(wire_d37_67),.data_out(wire_d37_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803769(.data_in(wire_d37_68),.data_out(wire_d37_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803770(.data_in(wire_d37_69),.data_out(wire_d37_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803771(.data_in(wire_d37_70),.data_out(wire_d37_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803772(.data_in(wire_d37_71),.data_out(wire_d37_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803773(.data_in(wire_d37_72),.data_out(wire_d37_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803774(.data_in(wire_d37_73),.data_out(wire_d37_74),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803775(.data_in(wire_d37_74),.data_out(wire_d37_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803776(.data_in(wire_d37_75),.data_out(wire_d37_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803777(.data_in(wire_d37_76),.data_out(wire_d37_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803778(.data_in(wire_d37_77),.data_out(wire_d37_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803779(.data_in(wire_d37_78),.data_out(d_out37),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance390380(.data_in(d_in38),.data_out(wire_d38_0),.clk(clk),.rst(rst));            //channel 39
	decoder_top #(.WIDTH(WIDTH)) decoder_instance390381(.data_in(wire_d38_0),.data_out(wire_d38_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance390382(.data_in(wire_d38_1),.data_out(wire_d38_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance390383(.data_in(wire_d38_2),.data_out(wire_d38_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance390384(.data_in(wire_d38_3),.data_out(wire_d38_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance390385(.data_in(wire_d38_4),.data_out(wire_d38_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance390386(.data_in(wire_d38_5),.data_out(wire_d38_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance390387(.data_in(wire_d38_6),.data_out(wire_d38_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance390388(.data_in(wire_d38_7),.data_out(wire_d38_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance390389(.data_in(wire_d38_8),.data_out(wire_d38_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903810(.data_in(wire_d38_9),.data_out(wire_d38_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903811(.data_in(wire_d38_10),.data_out(wire_d38_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903812(.data_in(wire_d38_11),.data_out(wire_d38_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903813(.data_in(wire_d38_12),.data_out(wire_d38_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903814(.data_in(wire_d38_13),.data_out(wire_d38_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903815(.data_in(wire_d38_14),.data_out(wire_d38_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903816(.data_in(wire_d38_15),.data_out(wire_d38_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903817(.data_in(wire_d38_16),.data_out(wire_d38_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903818(.data_in(wire_d38_17),.data_out(wire_d38_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903819(.data_in(wire_d38_18),.data_out(wire_d38_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903820(.data_in(wire_d38_19),.data_out(wire_d38_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903821(.data_in(wire_d38_20),.data_out(wire_d38_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903822(.data_in(wire_d38_21),.data_out(wire_d38_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903823(.data_in(wire_d38_22),.data_out(wire_d38_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903824(.data_in(wire_d38_23),.data_out(wire_d38_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903825(.data_in(wire_d38_24),.data_out(wire_d38_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903826(.data_in(wire_d38_25),.data_out(wire_d38_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903827(.data_in(wire_d38_26),.data_out(wire_d38_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903828(.data_in(wire_d38_27),.data_out(wire_d38_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903829(.data_in(wire_d38_28),.data_out(wire_d38_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903830(.data_in(wire_d38_29),.data_out(wire_d38_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903831(.data_in(wire_d38_30),.data_out(wire_d38_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903832(.data_in(wire_d38_31),.data_out(wire_d38_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903833(.data_in(wire_d38_32),.data_out(wire_d38_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903834(.data_in(wire_d38_33),.data_out(wire_d38_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903835(.data_in(wire_d38_34),.data_out(wire_d38_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903836(.data_in(wire_d38_35),.data_out(wire_d38_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903837(.data_in(wire_d38_36),.data_out(wire_d38_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903838(.data_in(wire_d38_37),.data_out(wire_d38_38),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903839(.data_in(wire_d38_38),.data_out(wire_d38_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903840(.data_in(wire_d38_39),.data_out(wire_d38_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903841(.data_in(wire_d38_40),.data_out(wire_d38_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903842(.data_in(wire_d38_41),.data_out(wire_d38_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903843(.data_in(wire_d38_42),.data_out(wire_d38_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903844(.data_in(wire_d38_43),.data_out(wire_d38_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903845(.data_in(wire_d38_44),.data_out(wire_d38_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903846(.data_in(wire_d38_45),.data_out(wire_d38_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903847(.data_in(wire_d38_46),.data_out(wire_d38_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903848(.data_in(wire_d38_47),.data_out(wire_d38_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903849(.data_in(wire_d38_48),.data_out(wire_d38_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903850(.data_in(wire_d38_49),.data_out(wire_d38_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903851(.data_in(wire_d38_50),.data_out(wire_d38_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903852(.data_in(wire_d38_51),.data_out(wire_d38_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903853(.data_in(wire_d38_52),.data_out(wire_d38_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903854(.data_in(wire_d38_53),.data_out(wire_d38_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903855(.data_in(wire_d38_54),.data_out(wire_d38_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903856(.data_in(wire_d38_55),.data_out(wire_d38_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903857(.data_in(wire_d38_56),.data_out(wire_d38_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903858(.data_in(wire_d38_57),.data_out(wire_d38_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903859(.data_in(wire_d38_58),.data_out(wire_d38_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903860(.data_in(wire_d38_59),.data_out(wire_d38_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903861(.data_in(wire_d38_60),.data_out(wire_d38_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903862(.data_in(wire_d38_61),.data_out(wire_d38_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903863(.data_in(wire_d38_62),.data_out(wire_d38_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903864(.data_in(wire_d38_63),.data_out(wire_d38_64),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903865(.data_in(wire_d38_64),.data_out(wire_d38_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903866(.data_in(wire_d38_65),.data_out(wire_d38_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903867(.data_in(wire_d38_66),.data_out(wire_d38_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903868(.data_in(wire_d38_67),.data_out(wire_d38_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903869(.data_in(wire_d38_68),.data_out(wire_d38_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903870(.data_in(wire_d38_69),.data_out(wire_d38_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903871(.data_in(wire_d38_70),.data_out(wire_d38_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903872(.data_in(wire_d38_71),.data_out(wire_d38_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903873(.data_in(wire_d38_72),.data_out(wire_d38_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903874(.data_in(wire_d38_73),.data_out(wire_d38_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903875(.data_in(wire_d38_74),.data_out(wire_d38_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903876(.data_in(wire_d38_75),.data_out(wire_d38_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903877(.data_in(wire_d38_76),.data_out(wire_d38_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903878(.data_in(wire_d38_77),.data_out(wire_d38_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903879(.data_in(wire_d38_78),.data_out(d_out38),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance400390(.data_in(d_in39),.data_out(wire_d39_0),.clk(clk),.rst(rst));            //channel 40
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance400391(.data_in(wire_d39_0),.data_out(wire_d39_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance400392(.data_in(wire_d39_1),.data_out(wire_d39_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance400393(.data_in(wire_d39_2),.data_out(wire_d39_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance400394(.data_in(wire_d39_3),.data_out(wire_d39_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance400395(.data_in(wire_d39_4),.data_out(wire_d39_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance400396(.data_in(wire_d39_5),.data_out(wire_d39_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance400397(.data_in(wire_d39_6),.data_out(wire_d39_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance400398(.data_in(wire_d39_7),.data_out(wire_d39_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance400399(.data_in(wire_d39_8),.data_out(wire_d39_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003910(.data_in(wire_d39_9),.data_out(wire_d39_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003911(.data_in(wire_d39_10),.data_out(wire_d39_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003912(.data_in(wire_d39_11),.data_out(wire_d39_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003913(.data_in(wire_d39_12),.data_out(wire_d39_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003914(.data_in(wire_d39_13),.data_out(wire_d39_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003915(.data_in(wire_d39_14),.data_out(wire_d39_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003916(.data_in(wire_d39_15),.data_out(wire_d39_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003917(.data_in(wire_d39_16),.data_out(wire_d39_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003918(.data_in(wire_d39_17),.data_out(wire_d39_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003919(.data_in(wire_d39_18),.data_out(wire_d39_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003920(.data_in(wire_d39_19),.data_out(wire_d39_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003921(.data_in(wire_d39_20),.data_out(wire_d39_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003922(.data_in(wire_d39_21),.data_out(wire_d39_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003923(.data_in(wire_d39_22),.data_out(wire_d39_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003924(.data_in(wire_d39_23),.data_out(wire_d39_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003925(.data_in(wire_d39_24),.data_out(wire_d39_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003926(.data_in(wire_d39_25),.data_out(wire_d39_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003927(.data_in(wire_d39_26),.data_out(wire_d39_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003928(.data_in(wire_d39_27),.data_out(wire_d39_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003929(.data_in(wire_d39_28),.data_out(wire_d39_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003930(.data_in(wire_d39_29),.data_out(wire_d39_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003931(.data_in(wire_d39_30),.data_out(wire_d39_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003932(.data_in(wire_d39_31),.data_out(wire_d39_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003933(.data_in(wire_d39_32),.data_out(wire_d39_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003934(.data_in(wire_d39_33),.data_out(wire_d39_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003935(.data_in(wire_d39_34),.data_out(wire_d39_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003936(.data_in(wire_d39_35),.data_out(wire_d39_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003937(.data_in(wire_d39_36),.data_out(wire_d39_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003938(.data_in(wire_d39_37),.data_out(wire_d39_38),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003939(.data_in(wire_d39_38),.data_out(wire_d39_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003940(.data_in(wire_d39_39),.data_out(wire_d39_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003941(.data_in(wire_d39_40),.data_out(wire_d39_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003942(.data_in(wire_d39_41),.data_out(wire_d39_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003943(.data_in(wire_d39_42),.data_out(wire_d39_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003944(.data_in(wire_d39_43),.data_out(wire_d39_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003945(.data_in(wire_d39_44),.data_out(wire_d39_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003946(.data_in(wire_d39_45),.data_out(wire_d39_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003947(.data_in(wire_d39_46),.data_out(wire_d39_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003948(.data_in(wire_d39_47),.data_out(wire_d39_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003949(.data_in(wire_d39_48),.data_out(wire_d39_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003950(.data_in(wire_d39_49),.data_out(wire_d39_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003951(.data_in(wire_d39_50),.data_out(wire_d39_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003952(.data_in(wire_d39_51),.data_out(wire_d39_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003953(.data_in(wire_d39_52),.data_out(wire_d39_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003954(.data_in(wire_d39_53),.data_out(wire_d39_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003955(.data_in(wire_d39_54),.data_out(wire_d39_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003956(.data_in(wire_d39_55),.data_out(wire_d39_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003957(.data_in(wire_d39_56),.data_out(wire_d39_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003958(.data_in(wire_d39_57),.data_out(wire_d39_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003959(.data_in(wire_d39_58),.data_out(wire_d39_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003960(.data_in(wire_d39_59),.data_out(wire_d39_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003961(.data_in(wire_d39_60),.data_out(wire_d39_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003962(.data_in(wire_d39_61),.data_out(wire_d39_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003963(.data_in(wire_d39_62),.data_out(wire_d39_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003964(.data_in(wire_d39_63),.data_out(wire_d39_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003965(.data_in(wire_d39_64),.data_out(wire_d39_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003966(.data_in(wire_d39_65),.data_out(wire_d39_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003967(.data_in(wire_d39_66),.data_out(wire_d39_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003968(.data_in(wire_d39_67),.data_out(wire_d39_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003969(.data_in(wire_d39_68),.data_out(wire_d39_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003970(.data_in(wire_d39_69),.data_out(wire_d39_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003971(.data_in(wire_d39_70),.data_out(wire_d39_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003972(.data_in(wire_d39_71),.data_out(wire_d39_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003973(.data_in(wire_d39_72),.data_out(wire_d39_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003974(.data_in(wire_d39_73),.data_out(wire_d39_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003975(.data_in(wire_d39_74),.data_out(wire_d39_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003976(.data_in(wire_d39_75),.data_out(wire_d39_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003977(.data_in(wire_d39_76),.data_out(wire_d39_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003978(.data_in(wire_d39_77),.data_out(wire_d39_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003979(.data_in(wire_d39_78),.data_out(d_out39),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance410400(.data_in(d_in40),.data_out(wire_d40_0),.clk(clk),.rst(rst));            //channel 41
	decoder_top #(.WIDTH(WIDTH)) decoder_instance410401(.data_in(wire_d40_0),.data_out(wire_d40_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance410402(.data_in(wire_d40_1),.data_out(wire_d40_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance410403(.data_in(wire_d40_2),.data_out(wire_d40_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance410404(.data_in(wire_d40_3),.data_out(wire_d40_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance410405(.data_in(wire_d40_4),.data_out(wire_d40_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance410406(.data_in(wire_d40_5),.data_out(wire_d40_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance410407(.data_in(wire_d40_6),.data_out(wire_d40_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance410408(.data_in(wire_d40_7),.data_out(wire_d40_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance410409(.data_in(wire_d40_8),.data_out(wire_d40_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104010(.data_in(wire_d40_9),.data_out(wire_d40_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104011(.data_in(wire_d40_10),.data_out(wire_d40_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104012(.data_in(wire_d40_11),.data_out(wire_d40_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104013(.data_in(wire_d40_12),.data_out(wire_d40_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104014(.data_in(wire_d40_13),.data_out(wire_d40_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104015(.data_in(wire_d40_14),.data_out(wire_d40_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104016(.data_in(wire_d40_15),.data_out(wire_d40_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104017(.data_in(wire_d40_16),.data_out(wire_d40_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104018(.data_in(wire_d40_17),.data_out(wire_d40_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104019(.data_in(wire_d40_18),.data_out(wire_d40_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104020(.data_in(wire_d40_19),.data_out(wire_d40_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104021(.data_in(wire_d40_20),.data_out(wire_d40_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104022(.data_in(wire_d40_21),.data_out(wire_d40_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104023(.data_in(wire_d40_22),.data_out(wire_d40_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104024(.data_in(wire_d40_23),.data_out(wire_d40_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104025(.data_in(wire_d40_24),.data_out(wire_d40_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104026(.data_in(wire_d40_25),.data_out(wire_d40_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104027(.data_in(wire_d40_26),.data_out(wire_d40_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104028(.data_in(wire_d40_27),.data_out(wire_d40_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104029(.data_in(wire_d40_28),.data_out(wire_d40_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104030(.data_in(wire_d40_29),.data_out(wire_d40_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104031(.data_in(wire_d40_30),.data_out(wire_d40_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104032(.data_in(wire_d40_31),.data_out(wire_d40_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104033(.data_in(wire_d40_32),.data_out(wire_d40_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104034(.data_in(wire_d40_33),.data_out(wire_d40_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104035(.data_in(wire_d40_34),.data_out(wire_d40_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104036(.data_in(wire_d40_35),.data_out(wire_d40_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104037(.data_in(wire_d40_36),.data_out(wire_d40_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104038(.data_in(wire_d40_37),.data_out(wire_d40_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104039(.data_in(wire_d40_38),.data_out(wire_d40_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104040(.data_in(wire_d40_39),.data_out(wire_d40_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104041(.data_in(wire_d40_40),.data_out(wire_d40_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104042(.data_in(wire_d40_41),.data_out(wire_d40_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104043(.data_in(wire_d40_42),.data_out(wire_d40_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104044(.data_in(wire_d40_43),.data_out(wire_d40_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104045(.data_in(wire_d40_44),.data_out(wire_d40_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104046(.data_in(wire_d40_45),.data_out(wire_d40_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104047(.data_in(wire_d40_46),.data_out(wire_d40_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104048(.data_in(wire_d40_47),.data_out(wire_d40_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104049(.data_in(wire_d40_48),.data_out(wire_d40_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104050(.data_in(wire_d40_49),.data_out(wire_d40_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104051(.data_in(wire_d40_50),.data_out(wire_d40_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104052(.data_in(wire_d40_51),.data_out(wire_d40_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104053(.data_in(wire_d40_52),.data_out(wire_d40_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104054(.data_in(wire_d40_53),.data_out(wire_d40_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104055(.data_in(wire_d40_54),.data_out(wire_d40_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104056(.data_in(wire_d40_55),.data_out(wire_d40_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104057(.data_in(wire_d40_56),.data_out(wire_d40_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104058(.data_in(wire_d40_57),.data_out(wire_d40_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104059(.data_in(wire_d40_58),.data_out(wire_d40_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104060(.data_in(wire_d40_59),.data_out(wire_d40_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104061(.data_in(wire_d40_60),.data_out(wire_d40_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104062(.data_in(wire_d40_61),.data_out(wire_d40_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104063(.data_in(wire_d40_62),.data_out(wire_d40_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104064(.data_in(wire_d40_63),.data_out(wire_d40_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104065(.data_in(wire_d40_64),.data_out(wire_d40_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104066(.data_in(wire_d40_65),.data_out(wire_d40_66),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104067(.data_in(wire_d40_66),.data_out(wire_d40_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104068(.data_in(wire_d40_67),.data_out(wire_d40_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104069(.data_in(wire_d40_68),.data_out(wire_d40_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104070(.data_in(wire_d40_69),.data_out(wire_d40_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104071(.data_in(wire_d40_70),.data_out(wire_d40_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104072(.data_in(wire_d40_71),.data_out(wire_d40_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104073(.data_in(wire_d40_72),.data_out(wire_d40_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104074(.data_in(wire_d40_73),.data_out(wire_d40_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104075(.data_in(wire_d40_74),.data_out(wire_d40_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104076(.data_in(wire_d40_75),.data_out(wire_d40_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104077(.data_in(wire_d40_76),.data_out(wire_d40_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104078(.data_in(wire_d40_77),.data_out(wire_d40_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104079(.data_in(wire_d40_78),.data_out(d_out40),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance420410(.data_in(d_in41),.data_out(wire_d41_0),.clk(clk),.rst(rst));            //channel 42
	decoder_top #(.WIDTH(WIDTH)) decoder_instance420411(.data_in(wire_d41_0),.data_out(wire_d41_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance420412(.data_in(wire_d41_1),.data_out(wire_d41_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance420413(.data_in(wire_d41_2),.data_out(wire_d41_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance420414(.data_in(wire_d41_3),.data_out(wire_d41_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance420415(.data_in(wire_d41_4),.data_out(wire_d41_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance420416(.data_in(wire_d41_5),.data_out(wire_d41_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance420417(.data_in(wire_d41_6),.data_out(wire_d41_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance420418(.data_in(wire_d41_7),.data_out(wire_d41_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance420419(.data_in(wire_d41_8),.data_out(wire_d41_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204110(.data_in(wire_d41_9),.data_out(wire_d41_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204111(.data_in(wire_d41_10),.data_out(wire_d41_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204112(.data_in(wire_d41_11),.data_out(wire_d41_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204113(.data_in(wire_d41_12),.data_out(wire_d41_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204114(.data_in(wire_d41_13),.data_out(wire_d41_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204115(.data_in(wire_d41_14),.data_out(wire_d41_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204116(.data_in(wire_d41_15),.data_out(wire_d41_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204117(.data_in(wire_d41_16),.data_out(wire_d41_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204118(.data_in(wire_d41_17),.data_out(wire_d41_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204119(.data_in(wire_d41_18),.data_out(wire_d41_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204120(.data_in(wire_d41_19),.data_out(wire_d41_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204121(.data_in(wire_d41_20),.data_out(wire_d41_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204122(.data_in(wire_d41_21),.data_out(wire_d41_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204123(.data_in(wire_d41_22),.data_out(wire_d41_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204124(.data_in(wire_d41_23),.data_out(wire_d41_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204125(.data_in(wire_d41_24),.data_out(wire_d41_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204126(.data_in(wire_d41_25),.data_out(wire_d41_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204127(.data_in(wire_d41_26),.data_out(wire_d41_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204128(.data_in(wire_d41_27),.data_out(wire_d41_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204129(.data_in(wire_d41_28),.data_out(wire_d41_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204130(.data_in(wire_d41_29),.data_out(wire_d41_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204131(.data_in(wire_d41_30),.data_out(wire_d41_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204132(.data_in(wire_d41_31),.data_out(wire_d41_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204133(.data_in(wire_d41_32),.data_out(wire_d41_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204134(.data_in(wire_d41_33),.data_out(wire_d41_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204135(.data_in(wire_d41_34),.data_out(wire_d41_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204136(.data_in(wire_d41_35),.data_out(wire_d41_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204137(.data_in(wire_d41_36),.data_out(wire_d41_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204138(.data_in(wire_d41_37),.data_out(wire_d41_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204139(.data_in(wire_d41_38),.data_out(wire_d41_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204140(.data_in(wire_d41_39),.data_out(wire_d41_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204141(.data_in(wire_d41_40),.data_out(wire_d41_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204142(.data_in(wire_d41_41),.data_out(wire_d41_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204143(.data_in(wire_d41_42),.data_out(wire_d41_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204144(.data_in(wire_d41_43),.data_out(wire_d41_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204145(.data_in(wire_d41_44),.data_out(wire_d41_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204146(.data_in(wire_d41_45),.data_out(wire_d41_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204147(.data_in(wire_d41_46),.data_out(wire_d41_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204148(.data_in(wire_d41_47),.data_out(wire_d41_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204149(.data_in(wire_d41_48),.data_out(wire_d41_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204150(.data_in(wire_d41_49),.data_out(wire_d41_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204151(.data_in(wire_d41_50),.data_out(wire_d41_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204152(.data_in(wire_d41_51),.data_out(wire_d41_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204153(.data_in(wire_d41_52),.data_out(wire_d41_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204154(.data_in(wire_d41_53),.data_out(wire_d41_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204155(.data_in(wire_d41_54),.data_out(wire_d41_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204156(.data_in(wire_d41_55),.data_out(wire_d41_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204157(.data_in(wire_d41_56),.data_out(wire_d41_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204158(.data_in(wire_d41_57),.data_out(wire_d41_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204159(.data_in(wire_d41_58),.data_out(wire_d41_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204160(.data_in(wire_d41_59),.data_out(wire_d41_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204161(.data_in(wire_d41_60),.data_out(wire_d41_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204162(.data_in(wire_d41_61),.data_out(wire_d41_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204163(.data_in(wire_d41_62),.data_out(wire_d41_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204164(.data_in(wire_d41_63),.data_out(wire_d41_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204165(.data_in(wire_d41_64),.data_out(wire_d41_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204166(.data_in(wire_d41_65),.data_out(wire_d41_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204167(.data_in(wire_d41_66),.data_out(wire_d41_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204168(.data_in(wire_d41_67),.data_out(wire_d41_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204169(.data_in(wire_d41_68),.data_out(wire_d41_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204170(.data_in(wire_d41_69),.data_out(wire_d41_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204171(.data_in(wire_d41_70),.data_out(wire_d41_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204172(.data_in(wire_d41_71),.data_out(wire_d41_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204173(.data_in(wire_d41_72),.data_out(wire_d41_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204174(.data_in(wire_d41_73),.data_out(wire_d41_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204175(.data_in(wire_d41_74),.data_out(wire_d41_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204176(.data_in(wire_d41_75),.data_out(wire_d41_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204177(.data_in(wire_d41_76),.data_out(wire_d41_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204178(.data_in(wire_d41_77),.data_out(wire_d41_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204179(.data_in(wire_d41_78),.data_out(d_out41),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance430420(.data_in(d_in42),.data_out(wire_d42_0),.clk(clk),.rst(rst));            //channel 43
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance430421(.data_in(wire_d42_0),.data_out(wire_d42_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance430422(.data_in(wire_d42_1),.data_out(wire_d42_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance430423(.data_in(wire_d42_2),.data_out(wire_d42_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance430424(.data_in(wire_d42_3),.data_out(wire_d42_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance430425(.data_in(wire_d42_4),.data_out(wire_d42_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance430426(.data_in(wire_d42_5),.data_out(wire_d42_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance430427(.data_in(wire_d42_6),.data_out(wire_d42_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance430428(.data_in(wire_d42_7),.data_out(wire_d42_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance430429(.data_in(wire_d42_8),.data_out(wire_d42_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304210(.data_in(wire_d42_9),.data_out(wire_d42_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304211(.data_in(wire_d42_10),.data_out(wire_d42_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4304212(.data_in(wire_d42_11),.data_out(wire_d42_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304213(.data_in(wire_d42_12),.data_out(wire_d42_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4304214(.data_in(wire_d42_13),.data_out(wire_d42_14),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304215(.data_in(wire_d42_14),.data_out(wire_d42_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304216(.data_in(wire_d42_15),.data_out(wire_d42_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304217(.data_in(wire_d42_16),.data_out(wire_d42_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304218(.data_in(wire_d42_17),.data_out(wire_d42_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304219(.data_in(wire_d42_18),.data_out(wire_d42_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304220(.data_in(wire_d42_19),.data_out(wire_d42_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304221(.data_in(wire_d42_20),.data_out(wire_d42_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304222(.data_in(wire_d42_21),.data_out(wire_d42_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304223(.data_in(wire_d42_22),.data_out(wire_d42_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304224(.data_in(wire_d42_23),.data_out(wire_d42_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304225(.data_in(wire_d42_24),.data_out(wire_d42_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304226(.data_in(wire_d42_25),.data_out(wire_d42_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4304227(.data_in(wire_d42_26),.data_out(wire_d42_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304228(.data_in(wire_d42_27),.data_out(wire_d42_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4304229(.data_in(wire_d42_28),.data_out(wire_d42_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304230(.data_in(wire_d42_29),.data_out(wire_d42_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304231(.data_in(wire_d42_30),.data_out(wire_d42_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304232(.data_in(wire_d42_31),.data_out(wire_d42_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304233(.data_in(wire_d42_32),.data_out(wire_d42_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304234(.data_in(wire_d42_33),.data_out(wire_d42_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304235(.data_in(wire_d42_34),.data_out(wire_d42_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304236(.data_in(wire_d42_35),.data_out(wire_d42_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304237(.data_in(wire_d42_36),.data_out(wire_d42_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304238(.data_in(wire_d42_37),.data_out(wire_d42_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304239(.data_in(wire_d42_38),.data_out(wire_d42_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304240(.data_in(wire_d42_39),.data_out(wire_d42_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304241(.data_in(wire_d42_40),.data_out(wire_d42_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304242(.data_in(wire_d42_41),.data_out(wire_d42_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304243(.data_in(wire_d42_42),.data_out(wire_d42_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304244(.data_in(wire_d42_43),.data_out(wire_d42_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304245(.data_in(wire_d42_44),.data_out(wire_d42_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304246(.data_in(wire_d42_45),.data_out(wire_d42_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304247(.data_in(wire_d42_46),.data_out(wire_d42_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304248(.data_in(wire_d42_47),.data_out(wire_d42_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304249(.data_in(wire_d42_48),.data_out(wire_d42_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304250(.data_in(wire_d42_49),.data_out(wire_d42_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304251(.data_in(wire_d42_50),.data_out(wire_d42_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304252(.data_in(wire_d42_51),.data_out(wire_d42_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304253(.data_in(wire_d42_52),.data_out(wire_d42_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304254(.data_in(wire_d42_53),.data_out(wire_d42_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304255(.data_in(wire_d42_54),.data_out(wire_d42_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304256(.data_in(wire_d42_55),.data_out(wire_d42_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304257(.data_in(wire_d42_56),.data_out(wire_d42_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304258(.data_in(wire_d42_57),.data_out(wire_d42_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304259(.data_in(wire_d42_58),.data_out(wire_d42_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304260(.data_in(wire_d42_59),.data_out(wire_d42_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304261(.data_in(wire_d42_60),.data_out(wire_d42_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304262(.data_in(wire_d42_61),.data_out(wire_d42_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304263(.data_in(wire_d42_62),.data_out(wire_d42_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304264(.data_in(wire_d42_63),.data_out(wire_d42_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304265(.data_in(wire_d42_64),.data_out(wire_d42_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304266(.data_in(wire_d42_65),.data_out(wire_d42_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304267(.data_in(wire_d42_66),.data_out(wire_d42_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304268(.data_in(wire_d42_67),.data_out(wire_d42_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304269(.data_in(wire_d42_68),.data_out(wire_d42_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304270(.data_in(wire_d42_69),.data_out(wire_d42_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304271(.data_in(wire_d42_70),.data_out(wire_d42_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304272(.data_in(wire_d42_71),.data_out(wire_d42_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304273(.data_in(wire_d42_72),.data_out(wire_d42_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304274(.data_in(wire_d42_73),.data_out(wire_d42_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304275(.data_in(wire_d42_74),.data_out(wire_d42_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304276(.data_in(wire_d42_75),.data_out(wire_d42_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304277(.data_in(wire_d42_76),.data_out(wire_d42_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304278(.data_in(wire_d42_77),.data_out(wire_d42_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304279(.data_in(wire_d42_78),.data_out(d_out42),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance440430(.data_in(d_in43),.data_out(wire_d43_0),.clk(clk),.rst(rst));            //channel 44
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance440431(.data_in(wire_d43_0),.data_out(wire_d43_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance440432(.data_in(wire_d43_1),.data_out(wire_d43_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance440433(.data_in(wire_d43_2),.data_out(wire_d43_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance440434(.data_in(wire_d43_3),.data_out(wire_d43_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance440435(.data_in(wire_d43_4),.data_out(wire_d43_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance440436(.data_in(wire_d43_5),.data_out(wire_d43_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance440437(.data_in(wire_d43_6),.data_out(wire_d43_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance440438(.data_in(wire_d43_7),.data_out(wire_d43_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance440439(.data_in(wire_d43_8),.data_out(wire_d43_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404310(.data_in(wire_d43_9),.data_out(wire_d43_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404311(.data_in(wire_d43_10),.data_out(wire_d43_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404312(.data_in(wire_d43_11),.data_out(wire_d43_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404313(.data_in(wire_d43_12),.data_out(wire_d43_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404314(.data_in(wire_d43_13),.data_out(wire_d43_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404315(.data_in(wire_d43_14),.data_out(wire_d43_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404316(.data_in(wire_d43_15),.data_out(wire_d43_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404317(.data_in(wire_d43_16),.data_out(wire_d43_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404318(.data_in(wire_d43_17),.data_out(wire_d43_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404319(.data_in(wire_d43_18),.data_out(wire_d43_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404320(.data_in(wire_d43_19),.data_out(wire_d43_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404321(.data_in(wire_d43_20),.data_out(wire_d43_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404322(.data_in(wire_d43_21),.data_out(wire_d43_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404323(.data_in(wire_d43_22),.data_out(wire_d43_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404324(.data_in(wire_d43_23),.data_out(wire_d43_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404325(.data_in(wire_d43_24),.data_out(wire_d43_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404326(.data_in(wire_d43_25),.data_out(wire_d43_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404327(.data_in(wire_d43_26),.data_out(wire_d43_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404328(.data_in(wire_d43_27),.data_out(wire_d43_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404329(.data_in(wire_d43_28),.data_out(wire_d43_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404330(.data_in(wire_d43_29),.data_out(wire_d43_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404331(.data_in(wire_d43_30),.data_out(wire_d43_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404332(.data_in(wire_d43_31),.data_out(wire_d43_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404333(.data_in(wire_d43_32),.data_out(wire_d43_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404334(.data_in(wire_d43_33),.data_out(wire_d43_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404335(.data_in(wire_d43_34),.data_out(wire_d43_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404336(.data_in(wire_d43_35),.data_out(wire_d43_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404337(.data_in(wire_d43_36),.data_out(wire_d43_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404338(.data_in(wire_d43_37),.data_out(wire_d43_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404339(.data_in(wire_d43_38),.data_out(wire_d43_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404340(.data_in(wire_d43_39),.data_out(wire_d43_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404341(.data_in(wire_d43_40),.data_out(wire_d43_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404342(.data_in(wire_d43_41),.data_out(wire_d43_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404343(.data_in(wire_d43_42),.data_out(wire_d43_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404344(.data_in(wire_d43_43),.data_out(wire_d43_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404345(.data_in(wire_d43_44),.data_out(wire_d43_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404346(.data_in(wire_d43_45),.data_out(wire_d43_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404347(.data_in(wire_d43_46),.data_out(wire_d43_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404348(.data_in(wire_d43_47),.data_out(wire_d43_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404349(.data_in(wire_d43_48),.data_out(wire_d43_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404350(.data_in(wire_d43_49),.data_out(wire_d43_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404351(.data_in(wire_d43_50),.data_out(wire_d43_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404352(.data_in(wire_d43_51),.data_out(wire_d43_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404353(.data_in(wire_d43_52),.data_out(wire_d43_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404354(.data_in(wire_d43_53),.data_out(wire_d43_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404355(.data_in(wire_d43_54),.data_out(wire_d43_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404356(.data_in(wire_d43_55),.data_out(wire_d43_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404357(.data_in(wire_d43_56),.data_out(wire_d43_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404358(.data_in(wire_d43_57),.data_out(wire_d43_58),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404359(.data_in(wire_d43_58),.data_out(wire_d43_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404360(.data_in(wire_d43_59),.data_out(wire_d43_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404361(.data_in(wire_d43_60),.data_out(wire_d43_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404362(.data_in(wire_d43_61),.data_out(wire_d43_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404363(.data_in(wire_d43_62),.data_out(wire_d43_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404364(.data_in(wire_d43_63),.data_out(wire_d43_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404365(.data_in(wire_d43_64),.data_out(wire_d43_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404366(.data_in(wire_d43_65),.data_out(wire_d43_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404367(.data_in(wire_d43_66),.data_out(wire_d43_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404368(.data_in(wire_d43_67),.data_out(wire_d43_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404369(.data_in(wire_d43_68),.data_out(wire_d43_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404370(.data_in(wire_d43_69),.data_out(wire_d43_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404371(.data_in(wire_d43_70),.data_out(wire_d43_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404372(.data_in(wire_d43_71),.data_out(wire_d43_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404373(.data_in(wire_d43_72),.data_out(wire_d43_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404374(.data_in(wire_d43_73),.data_out(wire_d43_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404375(.data_in(wire_d43_74),.data_out(wire_d43_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404376(.data_in(wire_d43_75),.data_out(wire_d43_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404377(.data_in(wire_d43_76),.data_out(wire_d43_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404378(.data_in(wire_d43_77),.data_out(wire_d43_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404379(.data_in(wire_d43_78),.data_out(d_out43),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance450440(.data_in(d_in44),.data_out(wire_d44_0),.clk(clk),.rst(rst));            //channel 45
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance450441(.data_in(wire_d44_0),.data_out(wire_d44_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance450442(.data_in(wire_d44_1),.data_out(wire_d44_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance450443(.data_in(wire_d44_2),.data_out(wire_d44_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance450444(.data_in(wire_d44_3),.data_out(wire_d44_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance450445(.data_in(wire_d44_4),.data_out(wire_d44_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance450446(.data_in(wire_d44_5),.data_out(wire_d44_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance450447(.data_in(wire_d44_6),.data_out(wire_d44_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance450448(.data_in(wire_d44_7),.data_out(wire_d44_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance450449(.data_in(wire_d44_8),.data_out(wire_d44_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504410(.data_in(wire_d44_9),.data_out(wire_d44_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504411(.data_in(wire_d44_10),.data_out(wire_d44_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504412(.data_in(wire_d44_11),.data_out(wire_d44_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504413(.data_in(wire_d44_12),.data_out(wire_d44_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504414(.data_in(wire_d44_13),.data_out(wire_d44_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504415(.data_in(wire_d44_14),.data_out(wire_d44_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504416(.data_in(wire_d44_15),.data_out(wire_d44_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504417(.data_in(wire_d44_16),.data_out(wire_d44_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504418(.data_in(wire_d44_17),.data_out(wire_d44_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504419(.data_in(wire_d44_18),.data_out(wire_d44_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504420(.data_in(wire_d44_19),.data_out(wire_d44_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504421(.data_in(wire_d44_20),.data_out(wire_d44_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504422(.data_in(wire_d44_21),.data_out(wire_d44_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504423(.data_in(wire_d44_22),.data_out(wire_d44_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504424(.data_in(wire_d44_23),.data_out(wire_d44_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504425(.data_in(wire_d44_24),.data_out(wire_d44_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504426(.data_in(wire_d44_25),.data_out(wire_d44_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504427(.data_in(wire_d44_26),.data_out(wire_d44_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504428(.data_in(wire_d44_27),.data_out(wire_d44_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504429(.data_in(wire_d44_28),.data_out(wire_d44_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504430(.data_in(wire_d44_29),.data_out(wire_d44_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504431(.data_in(wire_d44_30),.data_out(wire_d44_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504432(.data_in(wire_d44_31),.data_out(wire_d44_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504433(.data_in(wire_d44_32),.data_out(wire_d44_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504434(.data_in(wire_d44_33),.data_out(wire_d44_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504435(.data_in(wire_d44_34),.data_out(wire_d44_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504436(.data_in(wire_d44_35),.data_out(wire_d44_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504437(.data_in(wire_d44_36),.data_out(wire_d44_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504438(.data_in(wire_d44_37),.data_out(wire_d44_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504439(.data_in(wire_d44_38),.data_out(wire_d44_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504440(.data_in(wire_d44_39),.data_out(wire_d44_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504441(.data_in(wire_d44_40),.data_out(wire_d44_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504442(.data_in(wire_d44_41),.data_out(wire_d44_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504443(.data_in(wire_d44_42),.data_out(wire_d44_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504444(.data_in(wire_d44_43),.data_out(wire_d44_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504445(.data_in(wire_d44_44),.data_out(wire_d44_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504446(.data_in(wire_d44_45),.data_out(wire_d44_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504447(.data_in(wire_d44_46),.data_out(wire_d44_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504448(.data_in(wire_d44_47),.data_out(wire_d44_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504449(.data_in(wire_d44_48),.data_out(wire_d44_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504450(.data_in(wire_d44_49),.data_out(wire_d44_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504451(.data_in(wire_d44_50),.data_out(wire_d44_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504452(.data_in(wire_d44_51),.data_out(wire_d44_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504453(.data_in(wire_d44_52),.data_out(wire_d44_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504454(.data_in(wire_d44_53),.data_out(wire_d44_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504455(.data_in(wire_d44_54),.data_out(wire_d44_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504456(.data_in(wire_d44_55),.data_out(wire_d44_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504457(.data_in(wire_d44_56),.data_out(wire_d44_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504458(.data_in(wire_d44_57),.data_out(wire_d44_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504459(.data_in(wire_d44_58),.data_out(wire_d44_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504460(.data_in(wire_d44_59),.data_out(wire_d44_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504461(.data_in(wire_d44_60),.data_out(wire_d44_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504462(.data_in(wire_d44_61),.data_out(wire_d44_62),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504463(.data_in(wire_d44_62),.data_out(wire_d44_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504464(.data_in(wire_d44_63),.data_out(wire_d44_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504465(.data_in(wire_d44_64),.data_out(wire_d44_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504466(.data_in(wire_d44_65),.data_out(wire_d44_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504467(.data_in(wire_d44_66),.data_out(wire_d44_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504468(.data_in(wire_d44_67),.data_out(wire_d44_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504469(.data_in(wire_d44_68),.data_out(wire_d44_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504470(.data_in(wire_d44_69),.data_out(wire_d44_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504471(.data_in(wire_d44_70),.data_out(wire_d44_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504472(.data_in(wire_d44_71),.data_out(wire_d44_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504473(.data_in(wire_d44_72),.data_out(wire_d44_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504474(.data_in(wire_d44_73),.data_out(wire_d44_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504475(.data_in(wire_d44_74),.data_out(wire_d44_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504476(.data_in(wire_d44_75),.data_out(wire_d44_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504477(.data_in(wire_d44_76),.data_out(wire_d44_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504478(.data_in(wire_d44_77),.data_out(wire_d44_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504479(.data_in(wire_d44_78),.data_out(d_out44),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance460450(.data_in(d_in45),.data_out(wire_d45_0),.clk(clk),.rst(rst));            //channel 46
	decoder_top #(.WIDTH(WIDTH)) decoder_instance460451(.data_in(wire_d45_0),.data_out(wire_d45_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance460452(.data_in(wire_d45_1),.data_out(wire_d45_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance460453(.data_in(wire_d45_2),.data_out(wire_d45_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance460454(.data_in(wire_d45_3),.data_out(wire_d45_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance460455(.data_in(wire_d45_4),.data_out(wire_d45_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance460456(.data_in(wire_d45_5),.data_out(wire_d45_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance460457(.data_in(wire_d45_6),.data_out(wire_d45_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance460458(.data_in(wire_d45_7),.data_out(wire_d45_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance460459(.data_in(wire_d45_8),.data_out(wire_d45_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604510(.data_in(wire_d45_9),.data_out(wire_d45_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604511(.data_in(wire_d45_10),.data_out(wire_d45_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604512(.data_in(wire_d45_11),.data_out(wire_d45_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604513(.data_in(wire_d45_12),.data_out(wire_d45_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604514(.data_in(wire_d45_13),.data_out(wire_d45_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604515(.data_in(wire_d45_14),.data_out(wire_d45_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604516(.data_in(wire_d45_15),.data_out(wire_d45_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604517(.data_in(wire_d45_16),.data_out(wire_d45_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604518(.data_in(wire_d45_17),.data_out(wire_d45_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604519(.data_in(wire_d45_18),.data_out(wire_d45_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604520(.data_in(wire_d45_19),.data_out(wire_d45_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604521(.data_in(wire_d45_20),.data_out(wire_d45_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604522(.data_in(wire_d45_21),.data_out(wire_d45_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604523(.data_in(wire_d45_22),.data_out(wire_d45_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604524(.data_in(wire_d45_23),.data_out(wire_d45_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604525(.data_in(wire_d45_24),.data_out(wire_d45_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604526(.data_in(wire_d45_25),.data_out(wire_d45_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604527(.data_in(wire_d45_26),.data_out(wire_d45_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604528(.data_in(wire_d45_27),.data_out(wire_d45_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604529(.data_in(wire_d45_28),.data_out(wire_d45_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604530(.data_in(wire_d45_29),.data_out(wire_d45_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604531(.data_in(wire_d45_30),.data_out(wire_d45_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604532(.data_in(wire_d45_31),.data_out(wire_d45_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604533(.data_in(wire_d45_32),.data_out(wire_d45_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604534(.data_in(wire_d45_33),.data_out(wire_d45_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604535(.data_in(wire_d45_34),.data_out(wire_d45_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604536(.data_in(wire_d45_35),.data_out(wire_d45_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604537(.data_in(wire_d45_36),.data_out(wire_d45_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604538(.data_in(wire_d45_37),.data_out(wire_d45_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604539(.data_in(wire_d45_38),.data_out(wire_d45_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604540(.data_in(wire_d45_39),.data_out(wire_d45_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604541(.data_in(wire_d45_40),.data_out(wire_d45_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604542(.data_in(wire_d45_41),.data_out(wire_d45_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604543(.data_in(wire_d45_42),.data_out(wire_d45_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604544(.data_in(wire_d45_43),.data_out(wire_d45_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604545(.data_in(wire_d45_44),.data_out(wire_d45_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604546(.data_in(wire_d45_45),.data_out(wire_d45_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604547(.data_in(wire_d45_46),.data_out(wire_d45_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604548(.data_in(wire_d45_47),.data_out(wire_d45_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604549(.data_in(wire_d45_48),.data_out(wire_d45_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604550(.data_in(wire_d45_49),.data_out(wire_d45_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604551(.data_in(wire_d45_50),.data_out(wire_d45_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604552(.data_in(wire_d45_51),.data_out(wire_d45_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604553(.data_in(wire_d45_52),.data_out(wire_d45_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604554(.data_in(wire_d45_53),.data_out(wire_d45_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604555(.data_in(wire_d45_54),.data_out(wire_d45_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604556(.data_in(wire_d45_55),.data_out(wire_d45_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604557(.data_in(wire_d45_56),.data_out(wire_d45_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604558(.data_in(wire_d45_57),.data_out(wire_d45_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604559(.data_in(wire_d45_58),.data_out(wire_d45_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604560(.data_in(wire_d45_59),.data_out(wire_d45_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604561(.data_in(wire_d45_60),.data_out(wire_d45_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604562(.data_in(wire_d45_61),.data_out(wire_d45_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604563(.data_in(wire_d45_62),.data_out(wire_d45_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604564(.data_in(wire_d45_63),.data_out(wire_d45_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604565(.data_in(wire_d45_64),.data_out(wire_d45_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604566(.data_in(wire_d45_65),.data_out(wire_d45_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604567(.data_in(wire_d45_66),.data_out(wire_d45_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604568(.data_in(wire_d45_67),.data_out(wire_d45_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604569(.data_in(wire_d45_68),.data_out(wire_d45_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604570(.data_in(wire_d45_69),.data_out(wire_d45_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604571(.data_in(wire_d45_70),.data_out(wire_d45_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604572(.data_in(wire_d45_71),.data_out(wire_d45_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604573(.data_in(wire_d45_72),.data_out(wire_d45_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604574(.data_in(wire_d45_73),.data_out(wire_d45_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604575(.data_in(wire_d45_74),.data_out(wire_d45_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604576(.data_in(wire_d45_75),.data_out(wire_d45_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604577(.data_in(wire_d45_76),.data_out(wire_d45_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604578(.data_in(wire_d45_77),.data_out(wire_d45_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604579(.data_in(wire_d45_78),.data_out(d_out45),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance470460(.data_in(d_in46),.data_out(wire_d46_0),.clk(clk),.rst(rst));            //channel 47
	decoder_top #(.WIDTH(WIDTH)) decoder_instance470461(.data_in(wire_d46_0),.data_out(wire_d46_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance470462(.data_in(wire_d46_1),.data_out(wire_d46_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance470463(.data_in(wire_d46_2),.data_out(wire_d46_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance470464(.data_in(wire_d46_3),.data_out(wire_d46_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance470465(.data_in(wire_d46_4),.data_out(wire_d46_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance470466(.data_in(wire_d46_5),.data_out(wire_d46_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance470467(.data_in(wire_d46_6),.data_out(wire_d46_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance470468(.data_in(wire_d46_7),.data_out(wire_d46_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance470469(.data_in(wire_d46_8),.data_out(wire_d46_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704610(.data_in(wire_d46_9),.data_out(wire_d46_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704611(.data_in(wire_d46_10),.data_out(wire_d46_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704612(.data_in(wire_d46_11),.data_out(wire_d46_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704613(.data_in(wire_d46_12),.data_out(wire_d46_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704614(.data_in(wire_d46_13),.data_out(wire_d46_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704615(.data_in(wire_d46_14),.data_out(wire_d46_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704616(.data_in(wire_d46_15),.data_out(wire_d46_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704617(.data_in(wire_d46_16),.data_out(wire_d46_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704618(.data_in(wire_d46_17),.data_out(wire_d46_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704619(.data_in(wire_d46_18),.data_out(wire_d46_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704620(.data_in(wire_d46_19),.data_out(wire_d46_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704621(.data_in(wire_d46_20),.data_out(wire_d46_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704622(.data_in(wire_d46_21),.data_out(wire_d46_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704623(.data_in(wire_d46_22),.data_out(wire_d46_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704624(.data_in(wire_d46_23),.data_out(wire_d46_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704625(.data_in(wire_d46_24),.data_out(wire_d46_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704626(.data_in(wire_d46_25),.data_out(wire_d46_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704627(.data_in(wire_d46_26),.data_out(wire_d46_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704628(.data_in(wire_d46_27),.data_out(wire_d46_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704629(.data_in(wire_d46_28),.data_out(wire_d46_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704630(.data_in(wire_d46_29),.data_out(wire_d46_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704631(.data_in(wire_d46_30),.data_out(wire_d46_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704632(.data_in(wire_d46_31),.data_out(wire_d46_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704633(.data_in(wire_d46_32),.data_out(wire_d46_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704634(.data_in(wire_d46_33),.data_out(wire_d46_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704635(.data_in(wire_d46_34),.data_out(wire_d46_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704636(.data_in(wire_d46_35),.data_out(wire_d46_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704637(.data_in(wire_d46_36),.data_out(wire_d46_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704638(.data_in(wire_d46_37),.data_out(wire_d46_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704639(.data_in(wire_d46_38),.data_out(wire_d46_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704640(.data_in(wire_d46_39),.data_out(wire_d46_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704641(.data_in(wire_d46_40),.data_out(wire_d46_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704642(.data_in(wire_d46_41),.data_out(wire_d46_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704643(.data_in(wire_d46_42),.data_out(wire_d46_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704644(.data_in(wire_d46_43),.data_out(wire_d46_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704645(.data_in(wire_d46_44),.data_out(wire_d46_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704646(.data_in(wire_d46_45),.data_out(wire_d46_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704647(.data_in(wire_d46_46),.data_out(wire_d46_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704648(.data_in(wire_d46_47),.data_out(wire_d46_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704649(.data_in(wire_d46_48),.data_out(wire_d46_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704650(.data_in(wire_d46_49),.data_out(wire_d46_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704651(.data_in(wire_d46_50),.data_out(wire_d46_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704652(.data_in(wire_d46_51),.data_out(wire_d46_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704653(.data_in(wire_d46_52),.data_out(wire_d46_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704654(.data_in(wire_d46_53),.data_out(wire_d46_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704655(.data_in(wire_d46_54),.data_out(wire_d46_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704656(.data_in(wire_d46_55),.data_out(wire_d46_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704657(.data_in(wire_d46_56),.data_out(wire_d46_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704658(.data_in(wire_d46_57),.data_out(wire_d46_58),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704659(.data_in(wire_d46_58),.data_out(wire_d46_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704660(.data_in(wire_d46_59),.data_out(wire_d46_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704661(.data_in(wire_d46_60),.data_out(wire_d46_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704662(.data_in(wire_d46_61),.data_out(wire_d46_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704663(.data_in(wire_d46_62),.data_out(wire_d46_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704664(.data_in(wire_d46_63),.data_out(wire_d46_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704665(.data_in(wire_d46_64),.data_out(wire_d46_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704666(.data_in(wire_d46_65),.data_out(wire_d46_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704667(.data_in(wire_d46_66),.data_out(wire_d46_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704668(.data_in(wire_d46_67),.data_out(wire_d46_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704669(.data_in(wire_d46_68),.data_out(wire_d46_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704670(.data_in(wire_d46_69),.data_out(wire_d46_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704671(.data_in(wire_d46_70),.data_out(wire_d46_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704672(.data_in(wire_d46_71),.data_out(wire_d46_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704673(.data_in(wire_d46_72),.data_out(wire_d46_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704674(.data_in(wire_d46_73),.data_out(wire_d46_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704675(.data_in(wire_d46_74),.data_out(wire_d46_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704676(.data_in(wire_d46_75),.data_out(wire_d46_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704677(.data_in(wire_d46_76),.data_out(wire_d46_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704678(.data_in(wire_d46_77),.data_out(wire_d46_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704679(.data_in(wire_d46_78),.data_out(d_out46),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance480470(.data_in(d_in47),.data_out(wire_d47_0),.clk(clk),.rst(rst));            //channel 48
	invertion #(.WIDTH(WIDTH)) invertion_instance480471(.data_in(wire_d47_0),.data_out(wire_d47_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance480472(.data_in(wire_d47_1),.data_out(wire_d47_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance480473(.data_in(wire_d47_2),.data_out(wire_d47_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance480474(.data_in(wire_d47_3),.data_out(wire_d47_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance480475(.data_in(wire_d47_4),.data_out(wire_d47_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance480476(.data_in(wire_d47_5),.data_out(wire_d47_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance480477(.data_in(wire_d47_6),.data_out(wire_d47_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance480478(.data_in(wire_d47_7),.data_out(wire_d47_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance480479(.data_in(wire_d47_8),.data_out(wire_d47_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804710(.data_in(wire_d47_9),.data_out(wire_d47_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804711(.data_in(wire_d47_10),.data_out(wire_d47_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804712(.data_in(wire_d47_11),.data_out(wire_d47_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804713(.data_in(wire_d47_12),.data_out(wire_d47_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804714(.data_in(wire_d47_13),.data_out(wire_d47_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804715(.data_in(wire_d47_14),.data_out(wire_d47_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804716(.data_in(wire_d47_15),.data_out(wire_d47_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804717(.data_in(wire_d47_16),.data_out(wire_d47_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804718(.data_in(wire_d47_17),.data_out(wire_d47_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804719(.data_in(wire_d47_18),.data_out(wire_d47_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804720(.data_in(wire_d47_19),.data_out(wire_d47_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804721(.data_in(wire_d47_20),.data_out(wire_d47_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804722(.data_in(wire_d47_21),.data_out(wire_d47_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804723(.data_in(wire_d47_22),.data_out(wire_d47_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804724(.data_in(wire_d47_23),.data_out(wire_d47_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804725(.data_in(wire_d47_24),.data_out(wire_d47_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804726(.data_in(wire_d47_25),.data_out(wire_d47_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804727(.data_in(wire_d47_26),.data_out(wire_d47_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804728(.data_in(wire_d47_27),.data_out(wire_d47_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804729(.data_in(wire_d47_28),.data_out(wire_d47_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804730(.data_in(wire_d47_29),.data_out(wire_d47_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804731(.data_in(wire_d47_30),.data_out(wire_d47_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804732(.data_in(wire_d47_31),.data_out(wire_d47_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804733(.data_in(wire_d47_32),.data_out(wire_d47_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804734(.data_in(wire_d47_33),.data_out(wire_d47_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804735(.data_in(wire_d47_34),.data_out(wire_d47_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804736(.data_in(wire_d47_35),.data_out(wire_d47_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804737(.data_in(wire_d47_36),.data_out(wire_d47_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804738(.data_in(wire_d47_37),.data_out(wire_d47_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804739(.data_in(wire_d47_38),.data_out(wire_d47_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804740(.data_in(wire_d47_39),.data_out(wire_d47_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804741(.data_in(wire_d47_40),.data_out(wire_d47_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804742(.data_in(wire_d47_41),.data_out(wire_d47_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804743(.data_in(wire_d47_42),.data_out(wire_d47_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804744(.data_in(wire_d47_43),.data_out(wire_d47_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804745(.data_in(wire_d47_44),.data_out(wire_d47_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804746(.data_in(wire_d47_45),.data_out(wire_d47_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804747(.data_in(wire_d47_46),.data_out(wire_d47_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804748(.data_in(wire_d47_47),.data_out(wire_d47_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804749(.data_in(wire_d47_48),.data_out(wire_d47_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804750(.data_in(wire_d47_49),.data_out(wire_d47_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804751(.data_in(wire_d47_50),.data_out(wire_d47_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804752(.data_in(wire_d47_51),.data_out(wire_d47_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804753(.data_in(wire_d47_52),.data_out(wire_d47_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804754(.data_in(wire_d47_53),.data_out(wire_d47_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804755(.data_in(wire_d47_54),.data_out(wire_d47_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804756(.data_in(wire_d47_55),.data_out(wire_d47_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804757(.data_in(wire_d47_56),.data_out(wire_d47_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804758(.data_in(wire_d47_57),.data_out(wire_d47_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804759(.data_in(wire_d47_58),.data_out(wire_d47_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804760(.data_in(wire_d47_59),.data_out(wire_d47_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804761(.data_in(wire_d47_60),.data_out(wire_d47_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804762(.data_in(wire_d47_61),.data_out(wire_d47_62),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804763(.data_in(wire_d47_62),.data_out(wire_d47_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804764(.data_in(wire_d47_63),.data_out(wire_d47_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804765(.data_in(wire_d47_64),.data_out(wire_d47_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804766(.data_in(wire_d47_65),.data_out(wire_d47_66),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804767(.data_in(wire_d47_66),.data_out(wire_d47_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804768(.data_in(wire_d47_67),.data_out(wire_d47_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804769(.data_in(wire_d47_68),.data_out(wire_d47_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804770(.data_in(wire_d47_69),.data_out(wire_d47_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804771(.data_in(wire_d47_70),.data_out(wire_d47_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804772(.data_in(wire_d47_71),.data_out(wire_d47_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804773(.data_in(wire_d47_72),.data_out(wire_d47_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804774(.data_in(wire_d47_73),.data_out(wire_d47_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804775(.data_in(wire_d47_74),.data_out(wire_d47_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804776(.data_in(wire_d47_75),.data_out(wire_d47_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804777(.data_in(wire_d47_76),.data_out(wire_d47_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804778(.data_in(wire_d47_77),.data_out(wire_d47_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804779(.data_in(wire_d47_78),.data_out(d_out47),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance490480(.data_in(d_in48),.data_out(wire_d48_0),.clk(clk),.rst(rst));            //channel 49
	decoder_top #(.WIDTH(WIDTH)) decoder_instance490481(.data_in(wire_d48_0),.data_out(wire_d48_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance490482(.data_in(wire_d48_1),.data_out(wire_d48_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance490483(.data_in(wire_d48_2),.data_out(wire_d48_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance490484(.data_in(wire_d48_3),.data_out(wire_d48_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance490485(.data_in(wire_d48_4),.data_out(wire_d48_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance490486(.data_in(wire_d48_5),.data_out(wire_d48_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance490487(.data_in(wire_d48_6),.data_out(wire_d48_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance490488(.data_in(wire_d48_7),.data_out(wire_d48_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance490489(.data_in(wire_d48_8),.data_out(wire_d48_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904810(.data_in(wire_d48_9),.data_out(wire_d48_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904811(.data_in(wire_d48_10),.data_out(wire_d48_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904812(.data_in(wire_d48_11),.data_out(wire_d48_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904813(.data_in(wire_d48_12),.data_out(wire_d48_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904814(.data_in(wire_d48_13),.data_out(wire_d48_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904815(.data_in(wire_d48_14),.data_out(wire_d48_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904816(.data_in(wire_d48_15),.data_out(wire_d48_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904817(.data_in(wire_d48_16),.data_out(wire_d48_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904818(.data_in(wire_d48_17),.data_out(wire_d48_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904819(.data_in(wire_d48_18),.data_out(wire_d48_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904820(.data_in(wire_d48_19),.data_out(wire_d48_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904821(.data_in(wire_d48_20),.data_out(wire_d48_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904822(.data_in(wire_d48_21),.data_out(wire_d48_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904823(.data_in(wire_d48_22),.data_out(wire_d48_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904824(.data_in(wire_d48_23),.data_out(wire_d48_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904825(.data_in(wire_d48_24),.data_out(wire_d48_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904826(.data_in(wire_d48_25),.data_out(wire_d48_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904827(.data_in(wire_d48_26),.data_out(wire_d48_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904828(.data_in(wire_d48_27),.data_out(wire_d48_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904829(.data_in(wire_d48_28),.data_out(wire_d48_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904830(.data_in(wire_d48_29),.data_out(wire_d48_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904831(.data_in(wire_d48_30),.data_out(wire_d48_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904832(.data_in(wire_d48_31),.data_out(wire_d48_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904833(.data_in(wire_d48_32),.data_out(wire_d48_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904834(.data_in(wire_d48_33),.data_out(wire_d48_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904835(.data_in(wire_d48_34),.data_out(wire_d48_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904836(.data_in(wire_d48_35),.data_out(wire_d48_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904837(.data_in(wire_d48_36),.data_out(wire_d48_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904838(.data_in(wire_d48_37),.data_out(wire_d48_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904839(.data_in(wire_d48_38),.data_out(wire_d48_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904840(.data_in(wire_d48_39),.data_out(wire_d48_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904841(.data_in(wire_d48_40),.data_out(wire_d48_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904842(.data_in(wire_d48_41),.data_out(wire_d48_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904843(.data_in(wire_d48_42),.data_out(wire_d48_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904844(.data_in(wire_d48_43),.data_out(wire_d48_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904845(.data_in(wire_d48_44),.data_out(wire_d48_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904846(.data_in(wire_d48_45),.data_out(wire_d48_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904847(.data_in(wire_d48_46),.data_out(wire_d48_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904848(.data_in(wire_d48_47),.data_out(wire_d48_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904849(.data_in(wire_d48_48),.data_out(wire_d48_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904850(.data_in(wire_d48_49),.data_out(wire_d48_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904851(.data_in(wire_d48_50),.data_out(wire_d48_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904852(.data_in(wire_d48_51),.data_out(wire_d48_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904853(.data_in(wire_d48_52),.data_out(wire_d48_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904854(.data_in(wire_d48_53),.data_out(wire_d48_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904855(.data_in(wire_d48_54),.data_out(wire_d48_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904856(.data_in(wire_d48_55),.data_out(wire_d48_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904857(.data_in(wire_d48_56),.data_out(wire_d48_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904858(.data_in(wire_d48_57),.data_out(wire_d48_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904859(.data_in(wire_d48_58),.data_out(wire_d48_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904860(.data_in(wire_d48_59),.data_out(wire_d48_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904861(.data_in(wire_d48_60),.data_out(wire_d48_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904862(.data_in(wire_d48_61),.data_out(wire_d48_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904863(.data_in(wire_d48_62),.data_out(wire_d48_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904864(.data_in(wire_d48_63),.data_out(wire_d48_64),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904865(.data_in(wire_d48_64),.data_out(wire_d48_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904866(.data_in(wire_d48_65),.data_out(wire_d48_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904867(.data_in(wire_d48_66),.data_out(wire_d48_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904868(.data_in(wire_d48_67),.data_out(wire_d48_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904869(.data_in(wire_d48_68),.data_out(wire_d48_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904870(.data_in(wire_d48_69),.data_out(wire_d48_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904871(.data_in(wire_d48_70),.data_out(wire_d48_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904872(.data_in(wire_d48_71),.data_out(wire_d48_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904873(.data_in(wire_d48_72),.data_out(wire_d48_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904874(.data_in(wire_d48_73),.data_out(wire_d48_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904875(.data_in(wire_d48_74),.data_out(wire_d48_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904876(.data_in(wire_d48_75),.data_out(wire_d48_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904877(.data_in(wire_d48_76),.data_out(wire_d48_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904878(.data_in(wire_d48_77),.data_out(wire_d48_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904879(.data_in(wire_d48_78),.data_out(d_out48),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance500490(.data_in(d_in49),.data_out(wire_d49_0),.clk(clk),.rst(rst));            //channel 50
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance500491(.data_in(wire_d49_0),.data_out(wire_d49_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance500492(.data_in(wire_d49_1),.data_out(wire_d49_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance500493(.data_in(wire_d49_2),.data_out(wire_d49_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance500494(.data_in(wire_d49_3),.data_out(wire_d49_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance500495(.data_in(wire_d49_4),.data_out(wire_d49_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance500496(.data_in(wire_d49_5),.data_out(wire_d49_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance500497(.data_in(wire_d49_6),.data_out(wire_d49_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance500498(.data_in(wire_d49_7),.data_out(wire_d49_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance500499(.data_in(wire_d49_8),.data_out(wire_d49_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004910(.data_in(wire_d49_9),.data_out(wire_d49_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004911(.data_in(wire_d49_10),.data_out(wire_d49_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004912(.data_in(wire_d49_11),.data_out(wire_d49_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004913(.data_in(wire_d49_12),.data_out(wire_d49_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004914(.data_in(wire_d49_13),.data_out(wire_d49_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004915(.data_in(wire_d49_14),.data_out(wire_d49_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004916(.data_in(wire_d49_15),.data_out(wire_d49_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004917(.data_in(wire_d49_16),.data_out(wire_d49_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004918(.data_in(wire_d49_17),.data_out(wire_d49_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004919(.data_in(wire_d49_18),.data_out(wire_d49_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004920(.data_in(wire_d49_19),.data_out(wire_d49_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004921(.data_in(wire_d49_20),.data_out(wire_d49_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004922(.data_in(wire_d49_21),.data_out(wire_d49_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004923(.data_in(wire_d49_22),.data_out(wire_d49_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004924(.data_in(wire_d49_23),.data_out(wire_d49_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004925(.data_in(wire_d49_24),.data_out(wire_d49_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004926(.data_in(wire_d49_25),.data_out(wire_d49_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004927(.data_in(wire_d49_26),.data_out(wire_d49_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004928(.data_in(wire_d49_27),.data_out(wire_d49_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004929(.data_in(wire_d49_28),.data_out(wire_d49_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004930(.data_in(wire_d49_29),.data_out(wire_d49_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004931(.data_in(wire_d49_30),.data_out(wire_d49_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004932(.data_in(wire_d49_31),.data_out(wire_d49_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004933(.data_in(wire_d49_32),.data_out(wire_d49_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004934(.data_in(wire_d49_33),.data_out(wire_d49_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004935(.data_in(wire_d49_34),.data_out(wire_d49_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004936(.data_in(wire_d49_35),.data_out(wire_d49_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004937(.data_in(wire_d49_36),.data_out(wire_d49_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004938(.data_in(wire_d49_37),.data_out(wire_d49_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004939(.data_in(wire_d49_38),.data_out(wire_d49_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004940(.data_in(wire_d49_39),.data_out(wire_d49_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004941(.data_in(wire_d49_40),.data_out(wire_d49_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004942(.data_in(wire_d49_41),.data_out(wire_d49_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004943(.data_in(wire_d49_42),.data_out(wire_d49_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004944(.data_in(wire_d49_43),.data_out(wire_d49_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004945(.data_in(wire_d49_44),.data_out(wire_d49_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004946(.data_in(wire_d49_45),.data_out(wire_d49_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004947(.data_in(wire_d49_46),.data_out(wire_d49_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004948(.data_in(wire_d49_47),.data_out(wire_d49_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004949(.data_in(wire_d49_48),.data_out(wire_d49_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004950(.data_in(wire_d49_49),.data_out(wire_d49_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004951(.data_in(wire_d49_50),.data_out(wire_d49_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004952(.data_in(wire_d49_51),.data_out(wire_d49_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004953(.data_in(wire_d49_52),.data_out(wire_d49_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004954(.data_in(wire_d49_53),.data_out(wire_d49_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004955(.data_in(wire_d49_54),.data_out(wire_d49_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004956(.data_in(wire_d49_55),.data_out(wire_d49_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004957(.data_in(wire_d49_56),.data_out(wire_d49_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004958(.data_in(wire_d49_57),.data_out(wire_d49_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004959(.data_in(wire_d49_58),.data_out(wire_d49_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004960(.data_in(wire_d49_59),.data_out(wire_d49_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004961(.data_in(wire_d49_60),.data_out(wire_d49_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004962(.data_in(wire_d49_61),.data_out(wire_d49_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004963(.data_in(wire_d49_62),.data_out(wire_d49_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004964(.data_in(wire_d49_63),.data_out(wire_d49_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004965(.data_in(wire_d49_64),.data_out(wire_d49_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004966(.data_in(wire_d49_65),.data_out(wire_d49_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004967(.data_in(wire_d49_66),.data_out(wire_d49_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004968(.data_in(wire_d49_67),.data_out(wire_d49_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004969(.data_in(wire_d49_68),.data_out(wire_d49_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004970(.data_in(wire_d49_69),.data_out(wire_d49_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004971(.data_in(wire_d49_70),.data_out(wire_d49_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004972(.data_in(wire_d49_71),.data_out(wire_d49_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004973(.data_in(wire_d49_72),.data_out(wire_d49_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004974(.data_in(wire_d49_73),.data_out(wire_d49_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004975(.data_in(wire_d49_74),.data_out(wire_d49_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004976(.data_in(wire_d49_75),.data_out(wire_d49_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004977(.data_in(wire_d49_76),.data_out(wire_d49_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004978(.data_in(wire_d49_77),.data_out(wire_d49_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004979(.data_in(wire_d49_78),.data_out(d_out49),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance510500(.data_in(d_in50),.data_out(wire_d50_0),.clk(clk),.rst(rst));            //channel 51
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance510501(.data_in(wire_d50_0),.data_out(wire_d50_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance510502(.data_in(wire_d50_1),.data_out(wire_d50_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance510503(.data_in(wire_d50_2),.data_out(wire_d50_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance510504(.data_in(wire_d50_3),.data_out(wire_d50_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance510505(.data_in(wire_d50_4),.data_out(wire_d50_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance510506(.data_in(wire_d50_5),.data_out(wire_d50_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance510507(.data_in(wire_d50_6),.data_out(wire_d50_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance510508(.data_in(wire_d50_7),.data_out(wire_d50_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance510509(.data_in(wire_d50_8),.data_out(wire_d50_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105010(.data_in(wire_d50_9),.data_out(wire_d50_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105011(.data_in(wire_d50_10),.data_out(wire_d50_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105012(.data_in(wire_d50_11),.data_out(wire_d50_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105013(.data_in(wire_d50_12),.data_out(wire_d50_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105014(.data_in(wire_d50_13),.data_out(wire_d50_14),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105015(.data_in(wire_d50_14),.data_out(wire_d50_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105016(.data_in(wire_d50_15),.data_out(wire_d50_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105017(.data_in(wire_d50_16),.data_out(wire_d50_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105018(.data_in(wire_d50_17),.data_out(wire_d50_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105019(.data_in(wire_d50_18),.data_out(wire_d50_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105020(.data_in(wire_d50_19),.data_out(wire_d50_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105021(.data_in(wire_d50_20),.data_out(wire_d50_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105022(.data_in(wire_d50_21),.data_out(wire_d50_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105023(.data_in(wire_d50_22),.data_out(wire_d50_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105024(.data_in(wire_d50_23),.data_out(wire_d50_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105025(.data_in(wire_d50_24),.data_out(wire_d50_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105026(.data_in(wire_d50_25),.data_out(wire_d50_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105027(.data_in(wire_d50_26),.data_out(wire_d50_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105028(.data_in(wire_d50_27),.data_out(wire_d50_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105029(.data_in(wire_d50_28),.data_out(wire_d50_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105030(.data_in(wire_d50_29),.data_out(wire_d50_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105031(.data_in(wire_d50_30),.data_out(wire_d50_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105032(.data_in(wire_d50_31),.data_out(wire_d50_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105033(.data_in(wire_d50_32),.data_out(wire_d50_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105034(.data_in(wire_d50_33),.data_out(wire_d50_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105035(.data_in(wire_d50_34),.data_out(wire_d50_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105036(.data_in(wire_d50_35),.data_out(wire_d50_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105037(.data_in(wire_d50_36),.data_out(wire_d50_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105038(.data_in(wire_d50_37),.data_out(wire_d50_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105039(.data_in(wire_d50_38),.data_out(wire_d50_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105040(.data_in(wire_d50_39),.data_out(wire_d50_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105041(.data_in(wire_d50_40),.data_out(wire_d50_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105042(.data_in(wire_d50_41),.data_out(wire_d50_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105043(.data_in(wire_d50_42),.data_out(wire_d50_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105044(.data_in(wire_d50_43),.data_out(wire_d50_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105045(.data_in(wire_d50_44),.data_out(wire_d50_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105046(.data_in(wire_d50_45),.data_out(wire_d50_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105047(.data_in(wire_d50_46),.data_out(wire_d50_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105048(.data_in(wire_d50_47),.data_out(wire_d50_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105049(.data_in(wire_d50_48),.data_out(wire_d50_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105050(.data_in(wire_d50_49),.data_out(wire_d50_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105051(.data_in(wire_d50_50),.data_out(wire_d50_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105052(.data_in(wire_d50_51),.data_out(wire_d50_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105053(.data_in(wire_d50_52),.data_out(wire_d50_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105054(.data_in(wire_d50_53),.data_out(wire_d50_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105055(.data_in(wire_d50_54),.data_out(wire_d50_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105056(.data_in(wire_d50_55),.data_out(wire_d50_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105057(.data_in(wire_d50_56),.data_out(wire_d50_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105058(.data_in(wire_d50_57),.data_out(wire_d50_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105059(.data_in(wire_d50_58),.data_out(wire_d50_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105060(.data_in(wire_d50_59),.data_out(wire_d50_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105061(.data_in(wire_d50_60),.data_out(wire_d50_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105062(.data_in(wire_d50_61),.data_out(wire_d50_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105063(.data_in(wire_d50_62),.data_out(wire_d50_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105064(.data_in(wire_d50_63),.data_out(wire_d50_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105065(.data_in(wire_d50_64),.data_out(wire_d50_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105066(.data_in(wire_d50_65),.data_out(wire_d50_66),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105067(.data_in(wire_d50_66),.data_out(wire_d50_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105068(.data_in(wire_d50_67),.data_out(wire_d50_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105069(.data_in(wire_d50_68),.data_out(wire_d50_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105070(.data_in(wire_d50_69),.data_out(wire_d50_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105071(.data_in(wire_d50_70),.data_out(wire_d50_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105072(.data_in(wire_d50_71),.data_out(wire_d50_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105073(.data_in(wire_d50_72),.data_out(wire_d50_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105074(.data_in(wire_d50_73),.data_out(wire_d50_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105075(.data_in(wire_d50_74),.data_out(wire_d50_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105076(.data_in(wire_d50_75),.data_out(wire_d50_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105077(.data_in(wire_d50_76),.data_out(wire_d50_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105078(.data_in(wire_d50_77),.data_out(wire_d50_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105079(.data_in(wire_d50_78),.data_out(d_out50),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance520510(.data_in(d_in51),.data_out(wire_d51_0),.clk(clk),.rst(rst));            //channel 52
	register #(.WIDTH(WIDTH)) register_instance520511(.data_in(wire_d51_0),.data_out(wire_d51_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance520512(.data_in(wire_d51_1),.data_out(wire_d51_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance520513(.data_in(wire_d51_2),.data_out(wire_d51_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance520514(.data_in(wire_d51_3),.data_out(wire_d51_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance520515(.data_in(wire_d51_4),.data_out(wire_d51_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance520516(.data_in(wire_d51_5),.data_out(wire_d51_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance520517(.data_in(wire_d51_6),.data_out(wire_d51_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance520518(.data_in(wire_d51_7),.data_out(wire_d51_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance520519(.data_in(wire_d51_8),.data_out(wire_d51_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205110(.data_in(wire_d51_9),.data_out(wire_d51_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205111(.data_in(wire_d51_10),.data_out(wire_d51_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205112(.data_in(wire_d51_11),.data_out(wire_d51_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205113(.data_in(wire_d51_12),.data_out(wire_d51_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205114(.data_in(wire_d51_13),.data_out(wire_d51_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205115(.data_in(wire_d51_14),.data_out(wire_d51_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205116(.data_in(wire_d51_15),.data_out(wire_d51_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205117(.data_in(wire_d51_16),.data_out(wire_d51_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205118(.data_in(wire_d51_17),.data_out(wire_d51_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205119(.data_in(wire_d51_18),.data_out(wire_d51_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205120(.data_in(wire_d51_19),.data_out(wire_d51_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205121(.data_in(wire_d51_20),.data_out(wire_d51_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205122(.data_in(wire_d51_21),.data_out(wire_d51_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205123(.data_in(wire_d51_22),.data_out(wire_d51_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205124(.data_in(wire_d51_23),.data_out(wire_d51_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205125(.data_in(wire_d51_24),.data_out(wire_d51_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205126(.data_in(wire_d51_25),.data_out(wire_d51_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205127(.data_in(wire_d51_26),.data_out(wire_d51_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205128(.data_in(wire_d51_27),.data_out(wire_d51_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205129(.data_in(wire_d51_28),.data_out(wire_d51_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205130(.data_in(wire_d51_29),.data_out(wire_d51_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205131(.data_in(wire_d51_30),.data_out(wire_d51_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205132(.data_in(wire_d51_31),.data_out(wire_d51_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205133(.data_in(wire_d51_32),.data_out(wire_d51_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205134(.data_in(wire_d51_33),.data_out(wire_d51_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205135(.data_in(wire_d51_34),.data_out(wire_d51_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205136(.data_in(wire_d51_35),.data_out(wire_d51_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205137(.data_in(wire_d51_36),.data_out(wire_d51_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205138(.data_in(wire_d51_37),.data_out(wire_d51_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205139(.data_in(wire_d51_38),.data_out(wire_d51_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205140(.data_in(wire_d51_39),.data_out(wire_d51_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205141(.data_in(wire_d51_40),.data_out(wire_d51_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205142(.data_in(wire_d51_41),.data_out(wire_d51_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205143(.data_in(wire_d51_42),.data_out(wire_d51_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205144(.data_in(wire_d51_43),.data_out(wire_d51_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205145(.data_in(wire_d51_44),.data_out(wire_d51_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205146(.data_in(wire_d51_45),.data_out(wire_d51_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205147(.data_in(wire_d51_46),.data_out(wire_d51_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205148(.data_in(wire_d51_47),.data_out(wire_d51_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205149(.data_in(wire_d51_48),.data_out(wire_d51_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205150(.data_in(wire_d51_49),.data_out(wire_d51_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205151(.data_in(wire_d51_50),.data_out(wire_d51_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205152(.data_in(wire_d51_51),.data_out(wire_d51_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205153(.data_in(wire_d51_52),.data_out(wire_d51_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205154(.data_in(wire_d51_53),.data_out(wire_d51_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205155(.data_in(wire_d51_54),.data_out(wire_d51_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205156(.data_in(wire_d51_55),.data_out(wire_d51_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205157(.data_in(wire_d51_56),.data_out(wire_d51_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205158(.data_in(wire_d51_57),.data_out(wire_d51_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205159(.data_in(wire_d51_58),.data_out(wire_d51_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205160(.data_in(wire_d51_59),.data_out(wire_d51_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205161(.data_in(wire_d51_60),.data_out(wire_d51_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205162(.data_in(wire_d51_61),.data_out(wire_d51_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205163(.data_in(wire_d51_62),.data_out(wire_d51_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205164(.data_in(wire_d51_63),.data_out(wire_d51_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205165(.data_in(wire_d51_64),.data_out(wire_d51_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205166(.data_in(wire_d51_65),.data_out(wire_d51_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205167(.data_in(wire_d51_66),.data_out(wire_d51_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205168(.data_in(wire_d51_67),.data_out(wire_d51_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205169(.data_in(wire_d51_68),.data_out(wire_d51_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205170(.data_in(wire_d51_69),.data_out(wire_d51_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205171(.data_in(wire_d51_70),.data_out(wire_d51_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205172(.data_in(wire_d51_71),.data_out(wire_d51_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205173(.data_in(wire_d51_72),.data_out(wire_d51_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205174(.data_in(wire_d51_73),.data_out(wire_d51_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205175(.data_in(wire_d51_74),.data_out(wire_d51_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205176(.data_in(wire_d51_75),.data_out(wire_d51_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205177(.data_in(wire_d51_76),.data_out(wire_d51_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205178(.data_in(wire_d51_77),.data_out(wire_d51_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205179(.data_in(wire_d51_78),.data_out(d_out51),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance530520(.data_in(d_in52),.data_out(wire_d52_0),.clk(clk),.rst(rst));            //channel 53
	register #(.WIDTH(WIDTH)) register_instance530521(.data_in(wire_d52_0),.data_out(wire_d52_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance530522(.data_in(wire_d52_1),.data_out(wire_d52_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance530523(.data_in(wire_d52_2),.data_out(wire_d52_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance530524(.data_in(wire_d52_3),.data_out(wire_d52_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance530525(.data_in(wire_d52_4),.data_out(wire_d52_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance530526(.data_in(wire_d52_5),.data_out(wire_d52_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance530527(.data_in(wire_d52_6),.data_out(wire_d52_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance530528(.data_in(wire_d52_7),.data_out(wire_d52_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance530529(.data_in(wire_d52_8),.data_out(wire_d52_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305210(.data_in(wire_d52_9),.data_out(wire_d52_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305211(.data_in(wire_d52_10),.data_out(wire_d52_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305212(.data_in(wire_d52_11),.data_out(wire_d52_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305213(.data_in(wire_d52_12),.data_out(wire_d52_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305214(.data_in(wire_d52_13),.data_out(wire_d52_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305215(.data_in(wire_d52_14),.data_out(wire_d52_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305216(.data_in(wire_d52_15),.data_out(wire_d52_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305217(.data_in(wire_d52_16),.data_out(wire_d52_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305218(.data_in(wire_d52_17),.data_out(wire_d52_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305219(.data_in(wire_d52_18),.data_out(wire_d52_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305220(.data_in(wire_d52_19),.data_out(wire_d52_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305221(.data_in(wire_d52_20),.data_out(wire_d52_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305222(.data_in(wire_d52_21),.data_out(wire_d52_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305223(.data_in(wire_d52_22),.data_out(wire_d52_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305224(.data_in(wire_d52_23),.data_out(wire_d52_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305225(.data_in(wire_d52_24),.data_out(wire_d52_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305226(.data_in(wire_d52_25),.data_out(wire_d52_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305227(.data_in(wire_d52_26),.data_out(wire_d52_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305228(.data_in(wire_d52_27),.data_out(wire_d52_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305229(.data_in(wire_d52_28),.data_out(wire_d52_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305230(.data_in(wire_d52_29),.data_out(wire_d52_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305231(.data_in(wire_d52_30),.data_out(wire_d52_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305232(.data_in(wire_d52_31),.data_out(wire_d52_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305233(.data_in(wire_d52_32),.data_out(wire_d52_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305234(.data_in(wire_d52_33),.data_out(wire_d52_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305235(.data_in(wire_d52_34),.data_out(wire_d52_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305236(.data_in(wire_d52_35),.data_out(wire_d52_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305237(.data_in(wire_d52_36),.data_out(wire_d52_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305238(.data_in(wire_d52_37),.data_out(wire_d52_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305239(.data_in(wire_d52_38),.data_out(wire_d52_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305240(.data_in(wire_d52_39),.data_out(wire_d52_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305241(.data_in(wire_d52_40),.data_out(wire_d52_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305242(.data_in(wire_d52_41),.data_out(wire_d52_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305243(.data_in(wire_d52_42),.data_out(wire_d52_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305244(.data_in(wire_d52_43),.data_out(wire_d52_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305245(.data_in(wire_d52_44),.data_out(wire_d52_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305246(.data_in(wire_d52_45),.data_out(wire_d52_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305247(.data_in(wire_d52_46),.data_out(wire_d52_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305248(.data_in(wire_d52_47),.data_out(wire_d52_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305249(.data_in(wire_d52_48),.data_out(wire_d52_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305250(.data_in(wire_d52_49),.data_out(wire_d52_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305251(.data_in(wire_d52_50),.data_out(wire_d52_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305252(.data_in(wire_d52_51),.data_out(wire_d52_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305253(.data_in(wire_d52_52),.data_out(wire_d52_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305254(.data_in(wire_d52_53),.data_out(wire_d52_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305255(.data_in(wire_d52_54),.data_out(wire_d52_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305256(.data_in(wire_d52_55),.data_out(wire_d52_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305257(.data_in(wire_d52_56),.data_out(wire_d52_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305258(.data_in(wire_d52_57),.data_out(wire_d52_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305259(.data_in(wire_d52_58),.data_out(wire_d52_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305260(.data_in(wire_d52_59),.data_out(wire_d52_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305261(.data_in(wire_d52_60),.data_out(wire_d52_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305262(.data_in(wire_d52_61),.data_out(wire_d52_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305263(.data_in(wire_d52_62),.data_out(wire_d52_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305264(.data_in(wire_d52_63),.data_out(wire_d52_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305265(.data_in(wire_d52_64),.data_out(wire_d52_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305266(.data_in(wire_d52_65),.data_out(wire_d52_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305267(.data_in(wire_d52_66),.data_out(wire_d52_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305268(.data_in(wire_d52_67),.data_out(wire_d52_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305269(.data_in(wire_d52_68),.data_out(wire_d52_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305270(.data_in(wire_d52_69),.data_out(wire_d52_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305271(.data_in(wire_d52_70),.data_out(wire_d52_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305272(.data_in(wire_d52_71),.data_out(wire_d52_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305273(.data_in(wire_d52_72),.data_out(wire_d52_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305274(.data_in(wire_d52_73),.data_out(wire_d52_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305275(.data_in(wire_d52_74),.data_out(wire_d52_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305276(.data_in(wire_d52_75),.data_out(wire_d52_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305277(.data_in(wire_d52_76),.data_out(wire_d52_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305278(.data_in(wire_d52_77),.data_out(wire_d52_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305279(.data_in(wire_d52_78),.data_out(d_out52),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance540530(.data_in(d_in53),.data_out(wire_d53_0),.clk(clk),.rst(rst));            //channel 54
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance540531(.data_in(wire_d53_0),.data_out(wire_d53_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance540532(.data_in(wire_d53_1),.data_out(wire_d53_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance540533(.data_in(wire_d53_2),.data_out(wire_d53_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance540534(.data_in(wire_d53_3),.data_out(wire_d53_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance540535(.data_in(wire_d53_4),.data_out(wire_d53_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance540536(.data_in(wire_d53_5),.data_out(wire_d53_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance540537(.data_in(wire_d53_6),.data_out(wire_d53_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance540538(.data_in(wire_d53_7),.data_out(wire_d53_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance540539(.data_in(wire_d53_8),.data_out(wire_d53_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405310(.data_in(wire_d53_9),.data_out(wire_d53_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405311(.data_in(wire_d53_10),.data_out(wire_d53_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405312(.data_in(wire_d53_11),.data_out(wire_d53_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405313(.data_in(wire_d53_12),.data_out(wire_d53_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405314(.data_in(wire_d53_13),.data_out(wire_d53_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405315(.data_in(wire_d53_14),.data_out(wire_d53_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405316(.data_in(wire_d53_15),.data_out(wire_d53_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405317(.data_in(wire_d53_16),.data_out(wire_d53_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405318(.data_in(wire_d53_17),.data_out(wire_d53_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5405319(.data_in(wire_d53_18),.data_out(wire_d53_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405320(.data_in(wire_d53_19),.data_out(wire_d53_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405321(.data_in(wire_d53_20),.data_out(wire_d53_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405322(.data_in(wire_d53_21),.data_out(wire_d53_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405323(.data_in(wire_d53_22),.data_out(wire_d53_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405324(.data_in(wire_d53_23),.data_out(wire_d53_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405325(.data_in(wire_d53_24),.data_out(wire_d53_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405326(.data_in(wire_d53_25),.data_out(wire_d53_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405327(.data_in(wire_d53_26),.data_out(wire_d53_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405328(.data_in(wire_d53_27),.data_out(wire_d53_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405329(.data_in(wire_d53_28),.data_out(wire_d53_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405330(.data_in(wire_d53_29),.data_out(wire_d53_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405331(.data_in(wire_d53_30),.data_out(wire_d53_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405332(.data_in(wire_d53_31),.data_out(wire_d53_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405333(.data_in(wire_d53_32),.data_out(wire_d53_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5405334(.data_in(wire_d53_33),.data_out(wire_d53_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405335(.data_in(wire_d53_34),.data_out(wire_d53_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405336(.data_in(wire_d53_35),.data_out(wire_d53_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405337(.data_in(wire_d53_36),.data_out(wire_d53_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405338(.data_in(wire_d53_37),.data_out(wire_d53_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405339(.data_in(wire_d53_38),.data_out(wire_d53_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5405340(.data_in(wire_d53_39),.data_out(wire_d53_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405341(.data_in(wire_d53_40),.data_out(wire_d53_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405342(.data_in(wire_d53_41),.data_out(wire_d53_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405343(.data_in(wire_d53_42),.data_out(wire_d53_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405344(.data_in(wire_d53_43),.data_out(wire_d53_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405345(.data_in(wire_d53_44),.data_out(wire_d53_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405346(.data_in(wire_d53_45),.data_out(wire_d53_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405347(.data_in(wire_d53_46),.data_out(wire_d53_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405348(.data_in(wire_d53_47),.data_out(wire_d53_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405349(.data_in(wire_d53_48),.data_out(wire_d53_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405350(.data_in(wire_d53_49),.data_out(wire_d53_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405351(.data_in(wire_d53_50),.data_out(wire_d53_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405352(.data_in(wire_d53_51),.data_out(wire_d53_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405353(.data_in(wire_d53_52),.data_out(wire_d53_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5405354(.data_in(wire_d53_53),.data_out(wire_d53_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405355(.data_in(wire_d53_54),.data_out(wire_d53_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405356(.data_in(wire_d53_55),.data_out(wire_d53_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405357(.data_in(wire_d53_56),.data_out(wire_d53_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405358(.data_in(wire_d53_57),.data_out(wire_d53_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405359(.data_in(wire_d53_58),.data_out(wire_d53_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405360(.data_in(wire_d53_59),.data_out(wire_d53_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405361(.data_in(wire_d53_60),.data_out(wire_d53_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405362(.data_in(wire_d53_61),.data_out(wire_d53_62),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5405363(.data_in(wire_d53_62),.data_out(wire_d53_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405364(.data_in(wire_d53_63),.data_out(wire_d53_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405365(.data_in(wire_d53_64),.data_out(wire_d53_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405366(.data_in(wire_d53_65),.data_out(wire_d53_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405367(.data_in(wire_d53_66),.data_out(wire_d53_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405368(.data_in(wire_d53_67),.data_out(wire_d53_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405369(.data_in(wire_d53_68),.data_out(wire_d53_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405370(.data_in(wire_d53_69),.data_out(wire_d53_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405371(.data_in(wire_d53_70),.data_out(wire_d53_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405372(.data_in(wire_d53_71),.data_out(wire_d53_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405373(.data_in(wire_d53_72),.data_out(wire_d53_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405374(.data_in(wire_d53_73),.data_out(wire_d53_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405375(.data_in(wire_d53_74),.data_out(wire_d53_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405376(.data_in(wire_d53_75),.data_out(wire_d53_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405377(.data_in(wire_d53_76),.data_out(wire_d53_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405378(.data_in(wire_d53_77),.data_out(wire_d53_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405379(.data_in(wire_d53_78),.data_out(d_out53),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance550540(.data_in(d_in54),.data_out(wire_d54_0),.clk(clk),.rst(rst));            //channel 55
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance550541(.data_in(wire_d54_0),.data_out(wire_d54_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance550542(.data_in(wire_d54_1),.data_out(wire_d54_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance550543(.data_in(wire_d54_2),.data_out(wire_d54_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance550544(.data_in(wire_d54_3),.data_out(wire_d54_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance550545(.data_in(wire_d54_4),.data_out(wire_d54_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance550546(.data_in(wire_d54_5),.data_out(wire_d54_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance550547(.data_in(wire_d54_6),.data_out(wire_d54_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance550548(.data_in(wire_d54_7),.data_out(wire_d54_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance550549(.data_in(wire_d54_8),.data_out(wire_d54_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505410(.data_in(wire_d54_9),.data_out(wire_d54_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505411(.data_in(wire_d54_10),.data_out(wire_d54_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505412(.data_in(wire_d54_11),.data_out(wire_d54_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505413(.data_in(wire_d54_12),.data_out(wire_d54_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505414(.data_in(wire_d54_13),.data_out(wire_d54_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505415(.data_in(wire_d54_14),.data_out(wire_d54_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505416(.data_in(wire_d54_15),.data_out(wire_d54_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505417(.data_in(wire_d54_16),.data_out(wire_d54_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505418(.data_in(wire_d54_17),.data_out(wire_d54_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505419(.data_in(wire_d54_18),.data_out(wire_d54_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505420(.data_in(wire_d54_19),.data_out(wire_d54_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505421(.data_in(wire_d54_20),.data_out(wire_d54_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505422(.data_in(wire_d54_21),.data_out(wire_d54_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505423(.data_in(wire_d54_22),.data_out(wire_d54_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505424(.data_in(wire_d54_23),.data_out(wire_d54_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505425(.data_in(wire_d54_24),.data_out(wire_d54_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505426(.data_in(wire_d54_25),.data_out(wire_d54_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505427(.data_in(wire_d54_26),.data_out(wire_d54_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505428(.data_in(wire_d54_27),.data_out(wire_d54_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505429(.data_in(wire_d54_28),.data_out(wire_d54_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505430(.data_in(wire_d54_29),.data_out(wire_d54_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505431(.data_in(wire_d54_30),.data_out(wire_d54_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505432(.data_in(wire_d54_31),.data_out(wire_d54_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505433(.data_in(wire_d54_32),.data_out(wire_d54_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505434(.data_in(wire_d54_33),.data_out(wire_d54_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505435(.data_in(wire_d54_34),.data_out(wire_d54_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505436(.data_in(wire_d54_35),.data_out(wire_d54_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505437(.data_in(wire_d54_36),.data_out(wire_d54_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505438(.data_in(wire_d54_37),.data_out(wire_d54_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505439(.data_in(wire_d54_38),.data_out(wire_d54_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505440(.data_in(wire_d54_39),.data_out(wire_d54_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505441(.data_in(wire_d54_40),.data_out(wire_d54_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505442(.data_in(wire_d54_41),.data_out(wire_d54_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505443(.data_in(wire_d54_42),.data_out(wire_d54_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505444(.data_in(wire_d54_43),.data_out(wire_d54_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505445(.data_in(wire_d54_44),.data_out(wire_d54_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505446(.data_in(wire_d54_45),.data_out(wire_d54_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505447(.data_in(wire_d54_46),.data_out(wire_d54_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505448(.data_in(wire_d54_47),.data_out(wire_d54_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505449(.data_in(wire_d54_48),.data_out(wire_d54_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505450(.data_in(wire_d54_49),.data_out(wire_d54_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505451(.data_in(wire_d54_50),.data_out(wire_d54_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505452(.data_in(wire_d54_51),.data_out(wire_d54_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505453(.data_in(wire_d54_52),.data_out(wire_d54_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505454(.data_in(wire_d54_53),.data_out(wire_d54_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505455(.data_in(wire_d54_54),.data_out(wire_d54_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505456(.data_in(wire_d54_55),.data_out(wire_d54_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505457(.data_in(wire_d54_56),.data_out(wire_d54_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505458(.data_in(wire_d54_57),.data_out(wire_d54_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505459(.data_in(wire_d54_58),.data_out(wire_d54_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505460(.data_in(wire_d54_59),.data_out(wire_d54_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505461(.data_in(wire_d54_60),.data_out(wire_d54_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505462(.data_in(wire_d54_61),.data_out(wire_d54_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505463(.data_in(wire_d54_62),.data_out(wire_d54_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505464(.data_in(wire_d54_63),.data_out(wire_d54_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505465(.data_in(wire_d54_64),.data_out(wire_d54_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505466(.data_in(wire_d54_65),.data_out(wire_d54_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505467(.data_in(wire_d54_66),.data_out(wire_d54_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505468(.data_in(wire_d54_67),.data_out(wire_d54_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505469(.data_in(wire_d54_68),.data_out(wire_d54_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505470(.data_in(wire_d54_69),.data_out(wire_d54_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505471(.data_in(wire_d54_70),.data_out(wire_d54_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505472(.data_in(wire_d54_71),.data_out(wire_d54_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505473(.data_in(wire_d54_72),.data_out(wire_d54_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505474(.data_in(wire_d54_73),.data_out(wire_d54_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505475(.data_in(wire_d54_74),.data_out(wire_d54_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505476(.data_in(wire_d54_75),.data_out(wire_d54_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505477(.data_in(wire_d54_76),.data_out(wire_d54_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505478(.data_in(wire_d54_77),.data_out(wire_d54_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505479(.data_in(wire_d54_78),.data_out(d_out54),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance560550(.data_in(d_in55),.data_out(wire_d55_0),.clk(clk),.rst(rst));            //channel 56
	decoder_top #(.WIDTH(WIDTH)) decoder_instance560551(.data_in(wire_d55_0),.data_out(wire_d55_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance560552(.data_in(wire_d55_1),.data_out(wire_d55_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance560553(.data_in(wire_d55_2),.data_out(wire_d55_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance560554(.data_in(wire_d55_3),.data_out(wire_d55_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance560555(.data_in(wire_d55_4),.data_out(wire_d55_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance560556(.data_in(wire_d55_5),.data_out(wire_d55_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance560557(.data_in(wire_d55_6),.data_out(wire_d55_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance560558(.data_in(wire_d55_7),.data_out(wire_d55_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance560559(.data_in(wire_d55_8),.data_out(wire_d55_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605510(.data_in(wire_d55_9),.data_out(wire_d55_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605511(.data_in(wire_d55_10),.data_out(wire_d55_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605512(.data_in(wire_d55_11),.data_out(wire_d55_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605513(.data_in(wire_d55_12),.data_out(wire_d55_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605514(.data_in(wire_d55_13),.data_out(wire_d55_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605515(.data_in(wire_d55_14),.data_out(wire_d55_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605516(.data_in(wire_d55_15),.data_out(wire_d55_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605517(.data_in(wire_d55_16),.data_out(wire_d55_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605518(.data_in(wire_d55_17),.data_out(wire_d55_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605519(.data_in(wire_d55_18),.data_out(wire_d55_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605520(.data_in(wire_d55_19),.data_out(wire_d55_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605521(.data_in(wire_d55_20),.data_out(wire_d55_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605522(.data_in(wire_d55_21),.data_out(wire_d55_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605523(.data_in(wire_d55_22),.data_out(wire_d55_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605524(.data_in(wire_d55_23),.data_out(wire_d55_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605525(.data_in(wire_d55_24),.data_out(wire_d55_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605526(.data_in(wire_d55_25),.data_out(wire_d55_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605527(.data_in(wire_d55_26),.data_out(wire_d55_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605528(.data_in(wire_d55_27),.data_out(wire_d55_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605529(.data_in(wire_d55_28),.data_out(wire_d55_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605530(.data_in(wire_d55_29),.data_out(wire_d55_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605531(.data_in(wire_d55_30),.data_out(wire_d55_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605532(.data_in(wire_d55_31),.data_out(wire_d55_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605533(.data_in(wire_d55_32),.data_out(wire_d55_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605534(.data_in(wire_d55_33),.data_out(wire_d55_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605535(.data_in(wire_d55_34),.data_out(wire_d55_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605536(.data_in(wire_d55_35),.data_out(wire_d55_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605537(.data_in(wire_d55_36),.data_out(wire_d55_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605538(.data_in(wire_d55_37),.data_out(wire_d55_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605539(.data_in(wire_d55_38),.data_out(wire_d55_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605540(.data_in(wire_d55_39),.data_out(wire_d55_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605541(.data_in(wire_d55_40),.data_out(wire_d55_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605542(.data_in(wire_d55_41),.data_out(wire_d55_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605543(.data_in(wire_d55_42),.data_out(wire_d55_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605544(.data_in(wire_d55_43),.data_out(wire_d55_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605545(.data_in(wire_d55_44),.data_out(wire_d55_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605546(.data_in(wire_d55_45),.data_out(wire_d55_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605547(.data_in(wire_d55_46),.data_out(wire_d55_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605548(.data_in(wire_d55_47),.data_out(wire_d55_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605549(.data_in(wire_d55_48),.data_out(wire_d55_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605550(.data_in(wire_d55_49),.data_out(wire_d55_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605551(.data_in(wire_d55_50),.data_out(wire_d55_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605552(.data_in(wire_d55_51),.data_out(wire_d55_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605553(.data_in(wire_d55_52),.data_out(wire_d55_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605554(.data_in(wire_d55_53),.data_out(wire_d55_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605555(.data_in(wire_d55_54),.data_out(wire_d55_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605556(.data_in(wire_d55_55),.data_out(wire_d55_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605557(.data_in(wire_d55_56),.data_out(wire_d55_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605558(.data_in(wire_d55_57),.data_out(wire_d55_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605559(.data_in(wire_d55_58),.data_out(wire_d55_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605560(.data_in(wire_d55_59),.data_out(wire_d55_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605561(.data_in(wire_d55_60),.data_out(wire_d55_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605562(.data_in(wire_d55_61),.data_out(wire_d55_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605563(.data_in(wire_d55_62),.data_out(wire_d55_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605564(.data_in(wire_d55_63),.data_out(wire_d55_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605565(.data_in(wire_d55_64),.data_out(wire_d55_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605566(.data_in(wire_d55_65),.data_out(wire_d55_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605567(.data_in(wire_d55_66),.data_out(wire_d55_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605568(.data_in(wire_d55_67),.data_out(wire_d55_68),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605569(.data_in(wire_d55_68),.data_out(wire_d55_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605570(.data_in(wire_d55_69),.data_out(wire_d55_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605571(.data_in(wire_d55_70),.data_out(wire_d55_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605572(.data_in(wire_d55_71),.data_out(wire_d55_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605573(.data_in(wire_d55_72),.data_out(wire_d55_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605574(.data_in(wire_d55_73),.data_out(wire_d55_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605575(.data_in(wire_d55_74),.data_out(wire_d55_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605576(.data_in(wire_d55_75),.data_out(wire_d55_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605577(.data_in(wire_d55_76),.data_out(wire_d55_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605578(.data_in(wire_d55_77),.data_out(wire_d55_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605579(.data_in(wire_d55_78),.data_out(d_out55),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance570560(.data_in(d_in56),.data_out(wire_d56_0),.clk(clk),.rst(rst));            //channel 57
	register #(.WIDTH(WIDTH)) register_instance570561(.data_in(wire_d56_0),.data_out(wire_d56_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance570562(.data_in(wire_d56_1),.data_out(wire_d56_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance570563(.data_in(wire_d56_2),.data_out(wire_d56_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance570564(.data_in(wire_d56_3),.data_out(wire_d56_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance570565(.data_in(wire_d56_4),.data_out(wire_d56_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance570566(.data_in(wire_d56_5),.data_out(wire_d56_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance570567(.data_in(wire_d56_6),.data_out(wire_d56_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance570568(.data_in(wire_d56_7),.data_out(wire_d56_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance570569(.data_in(wire_d56_8),.data_out(wire_d56_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705610(.data_in(wire_d56_9),.data_out(wire_d56_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705611(.data_in(wire_d56_10),.data_out(wire_d56_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705612(.data_in(wire_d56_11),.data_out(wire_d56_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705613(.data_in(wire_d56_12),.data_out(wire_d56_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705614(.data_in(wire_d56_13),.data_out(wire_d56_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705615(.data_in(wire_d56_14),.data_out(wire_d56_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705616(.data_in(wire_d56_15),.data_out(wire_d56_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705617(.data_in(wire_d56_16),.data_out(wire_d56_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705618(.data_in(wire_d56_17),.data_out(wire_d56_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705619(.data_in(wire_d56_18),.data_out(wire_d56_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705620(.data_in(wire_d56_19),.data_out(wire_d56_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705621(.data_in(wire_d56_20),.data_out(wire_d56_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705622(.data_in(wire_d56_21),.data_out(wire_d56_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705623(.data_in(wire_d56_22),.data_out(wire_d56_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705624(.data_in(wire_d56_23),.data_out(wire_d56_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705625(.data_in(wire_d56_24),.data_out(wire_d56_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5705626(.data_in(wire_d56_25),.data_out(wire_d56_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705627(.data_in(wire_d56_26),.data_out(wire_d56_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705628(.data_in(wire_d56_27),.data_out(wire_d56_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705629(.data_in(wire_d56_28),.data_out(wire_d56_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5705630(.data_in(wire_d56_29),.data_out(wire_d56_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705631(.data_in(wire_d56_30),.data_out(wire_d56_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705632(.data_in(wire_d56_31),.data_out(wire_d56_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705633(.data_in(wire_d56_32),.data_out(wire_d56_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705634(.data_in(wire_d56_33),.data_out(wire_d56_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705635(.data_in(wire_d56_34),.data_out(wire_d56_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705636(.data_in(wire_d56_35),.data_out(wire_d56_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5705637(.data_in(wire_d56_36),.data_out(wire_d56_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705638(.data_in(wire_d56_37),.data_out(wire_d56_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705639(.data_in(wire_d56_38),.data_out(wire_d56_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705640(.data_in(wire_d56_39),.data_out(wire_d56_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705641(.data_in(wire_d56_40),.data_out(wire_d56_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705642(.data_in(wire_d56_41),.data_out(wire_d56_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705643(.data_in(wire_d56_42),.data_out(wire_d56_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5705644(.data_in(wire_d56_43),.data_out(wire_d56_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705645(.data_in(wire_d56_44),.data_out(wire_d56_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705646(.data_in(wire_d56_45),.data_out(wire_d56_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705647(.data_in(wire_d56_46),.data_out(wire_d56_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705648(.data_in(wire_d56_47),.data_out(wire_d56_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705649(.data_in(wire_d56_48),.data_out(wire_d56_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705650(.data_in(wire_d56_49),.data_out(wire_d56_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705651(.data_in(wire_d56_50),.data_out(wire_d56_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705652(.data_in(wire_d56_51),.data_out(wire_d56_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705653(.data_in(wire_d56_52),.data_out(wire_d56_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705654(.data_in(wire_d56_53),.data_out(wire_d56_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705655(.data_in(wire_d56_54),.data_out(wire_d56_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705656(.data_in(wire_d56_55),.data_out(wire_d56_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705657(.data_in(wire_d56_56),.data_out(wire_d56_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705658(.data_in(wire_d56_57),.data_out(wire_d56_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705659(.data_in(wire_d56_58),.data_out(wire_d56_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705660(.data_in(wire_d56_59),.data_out(wire_d56_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705661(.data_in(wire_d56_60),.data_out(wire_d56_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705662(.data_in(wire_d56_61),.data_out(wire_d56_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705663(.data_in(wire_d56_62),.data_out(wire_d56_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705664(.data_in(wire_d56_63),.data_out(wire_d56_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705665(.data_in(wire_d56_64),.data_out(wire_d56_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5705666(.data_in(wire_d56_65),.data_out(wire_d56_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705667(.data_in(wire_d56_66),.data_out(wire_d56_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705668(.data_in(wire_d56_67),.data_out(wire_d56_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705669(.data_in(wire_d56_68),.data_out(wire_d56_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705670(.data_in(wire_d56_69),.data_out(wire_d56_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705671(.data_in(wire_d56_70),.data_out(wire_d56_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705672(.data_in(wire_d56_71),.data_out(wire_d56_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705673(.data_in(wire_d56_72),.data_out(wire_d56_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705674(.data_in(wire_d56_73),.data_out(wire_d56_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705675(.data_in(wire_d56_74),.data_out(wire_d56_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705676(.data_in(wire_d56_75),.data_out(wire_d56_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705677(.data_in(wire_d56_76),.data_out(wire_d56_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705678(.data_in(wire_d56_77),.data_out(wire_d56_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705679(.data_in(wire_d56_78),.data_out(d_out56),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance580570(.data_in(d_in57),.data_out(wire_d57_0),.clk(clk),.rst(rst));            //channel 58
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance580571(.data_in(wire_d57_0),.data_out(wire_d57_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance580572(.data_in(wire_d57_1),.data_out(wire_d57_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance580573(.data_in(wire_d57_2),.data_out(wire_d57_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance580574(.data_in(wire_d57_3),.data_out(wire_d57_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance580575(.data_in(wire_d57_4),.data_out(wire_d57_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance580576(.data_in(wire_d57_5),.data_out(wire_d57_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance580577(.data_in(wire_d57_6),.data_out(wire_d57_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance580578(.data_in(wire_d57_7),.data_out(wire_d57_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance580579(.data_in(wire_d57_8),.data_out(wire_d57_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805710(.data_in(wire_d57_9),.data_out(wire_d57_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805711(.data_in(wire_d57_10),.data_out(wire_d57_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805712(.data_in(wire_d57_11),.data_out(wire_d57_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805713(.data_in(wire_d57_12),.data_out(wire_d57_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805714(.data_in(wire_d57_13),.data_out(wire_d57_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805715(.data_in(wire_d57_14),.data_out(wire_d57_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805716(.data_in(wire_d57_15),.data_out(wire_d57_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805717(.data_in(wire_d57_16),.data_out(wire_d57_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805718(.data_in(wire_d57_17),.data_out(wire_d57_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805719(.data_in(wire_d57_18),.data_out(wire_d57_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805720(.data_in(wire_d57_19),.data_out(wire_d57_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805721(.data_in(wire_d57_20),.data_out(wire_d57_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805722(.data_in(wire_d57_21),.data_out(wire_d57_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805723(.data_in(wire_d57_22),.data_out(wire_d57_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805724(.data_in(wire_d57_23),.data_out(wire_d57_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805725(.data_in(wire_d57_24),.data_out(wire_d57_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805726(.data_in(wire_d57_25),.data_out(wire_d57_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805727(.data_in(wire_d57_26),.data_out(wire_d57_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805728(.data_in(wire_d57_27),.data_out(wire_d57_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805729(.data_in(wire_d57_28),.data_out(wire_d57_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805730(.data_in(wire_d57_29),.data_out(wire_d57_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805731(.data_in(wire_d57_30),.data_out(wire_d57_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805732(.data_in(wire_d57_31),.data_out(wire_d57_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805733(.data_in(wire_d57_32),.data_out(wire_d57_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805734(.data_in(wire_d57_33),.data_out(wire_d57_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805735(.data_in(wire_d57_34),.data_out(wire_d57_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805736(.data_in(wire_d57_35),.data_out(wire_d57_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805737(.data_in(wire_d57_36),.data_out(wire_d57_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805738(.data_in(wire_d57_37),.data_out(wire_d57_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805739(.data_in(wire_d57_38),.data_out(wire_d57_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805740(.data_in(wire_d57_39),.data_out(wire_d57_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805741(.data_in(wire_d57_40),.data_out(wire_d57_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805742(.data_in(wire_d57_41),.data_out(wire_d57_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805743(.data_in(wire_d57_42),.data_out(wire_d57_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805744(.data_in(wire_d57_43),.data_out(wire_d57_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805745(.data_in(wire_d57_44),.data_out(wire_d57_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805746(.data_in(wire_d57_45),.data_out(wire_d57_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805747(.data_in(wire_d57_46),.data_out(wire_d57_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805748(.data_in(wire_d57_47),.data_out(wire_d57_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805749(.data_in(wire_d57_48),.data_out(wire_d57_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805750(.data_in(wire_d57_49),.data_out(wire_d57_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805751(.data_in(wire_d57_50),.data_out(wire_d57_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805752(.data_in(wire_d57_51),.data_out(wire_d57_52),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805753(.data_in(wire_d57_52),.data_out(wire_d57_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805754(.data_in(wire_d57_53),.data_out(wire_d57_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805755(.data_in(wire_d57_54),.data_out(wire_d57_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805756(.data_in(wire_d57_55),.data_out(wire_d57_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805757(.data_in(wire_d57_56),.data_out(wire_d57_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805758(.data_in(wire_d57_57),.data_out(wire_d57_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805759(.data_in(wire_d57_58),.data_out(wire_d57_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805760(.data_in(wire_d57_59),.data_out(wire_d57_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805761(.data_in(wire_d57_60),.data_out(wire_d57_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805762(.data_in(wire_d57_61),.data_out(wire_d57_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805763(.data_in(wire_d57_62),.data_out(wire_d57_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805764(.data_in(wire_d57_63),.data_out(wire_d57_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805765(.data_in(wire_d57_64),.data_out(wire_d57_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805766(.data_in(wire_d57_65),.data_out(wire_d57_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805767(.data_in(wire_d57_66),.data_out(wire_d57_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805768(.data_in(wire_d57_67),.data_out(wire_d57_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805769(.data_in(wire_d57_68),.data_out(wire_d57_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805770(.data_in(wire_d57_69),.data_out(wire_d57_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805771(.data_in(wire_d57_70),.data_out(wire_d57_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805772(.data_in(wire_d57_71),.data_out(wire_d57_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805773(.data_in(wire_d57_72),.data_out(wire_d57_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805774(.data_in(wire_d57_73),.data_out(wire_d57_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805775(.data_in(wire_d57_74),.data_out(wire_d57_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805776(.data_in(wire_d57_75),.data_out(wire_d57_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805777(.data_in(wire_d57_76),.data_out(wire_d57_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805778(.data_in(wire_d57_77),.data_out(wire_d57_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805779(.data_in(wire_d57_78),.data_out(d_out57),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance590580(.data_in(d_in58),.data_out(wire_d58_0),.clk(clk),.rst(rst));            //channel 59
	encoder #(.WIDTH(WIDTH)) encoder_instance590581(.data_in(wire_d58_0),.data_out(wire_d58_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance590582(.data_in(wire_d58_1),.data_out(wire_d58_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance590583(.data_in(wire_d58_2),.data_out(wire_d58_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance590584(.data_in(wire_d58_3),.data_out(wire_d58_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance590585(.data_in(wire_d58_4),.data_out(wire_d58_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance590586(.data_in(wire_d58_5),.data_out(wire_d58_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance590587(.data_in(wire_d58_6),.data_out(wire_d58_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance590588(.data_in(wire_d58_7),.data_out(wire_d58_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance590589(.data_in(wire_d58_8),.data_out(wire_d58_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905810(.data_in(wire_d58_9),.data_out(wire_d58_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905811(.data_in(wire_d58_10),.data_out(wire_d58_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905812(.data_in(wire_d58_11),.data_out(wire_d58_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905813(.data_in(wire_d58_12),.data_out(wire_d58_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905814(.data_in(wire_d58_13),.data_out(wire_d58_14),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905815(.data_in(wire_d58_14),.data_out(wire_d58_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905816(.data_in(wire_d58_15),.data_out(wire_d58_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905817(.data_in(wire_d58_16),.data_out(wire_d58_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905818(.data_in(wire_d58_17),.data_out(wire_d58_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905819(.data_in(wire_d58_18),.data_out(wire_d58_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905820(.data_in(wire_d58_19),.data_out(wire_d58_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905821(.data_in(wire_d58_20),.data_out(wire_d58_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905822(.data_in(wire_d58_21),.data_out(wire_d58_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905823(.data_in(wire_d58_22),.data_out(wire_d58_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905824(.data_in(wire_d58_23),.data_out(wire_d58_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905825(.data_in(wire_d58_24),.data_out(wire_d58_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905826(.data_in(wire_d58_25),.data_out(wire_d58_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905827(.data_in(wire_d58_26),.data_out(wire_d58_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905828(.data_in(wire_d58_27),.data_out(wire_d58_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905829(.data_in(wire_d58_28),.data_out(wire_d58_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905830(.data_in(wire_d58_29),.data_out(wire_d58_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905831(.data_in(wire_d58_30),.data_out(wire_d58_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905832(.data_in(wire_d58_31),.data_out(wire_d58_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905833(.data_in(wire_d58_32),.data_out(wire_d58_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905834(.data_in(wire_d58_33),.data_out(wire_d58_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905835(.data_in(wire_d58_34),.data_out(wire_d58_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905836(.data_in(wire_d58_35),.data_out(wire_d58_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905837(.data_in(wire_d58_36),.data_out(wire_d58_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905838(.data_in(wire_d58_37),.data_out(wire_d58_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905839(.data_in(wire_d58_38),.data_out(wire_d58_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905840(.data_in(wire_d58_39),.data_out(wire_d58_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905841(.data_in(wire_d58_40),.data_out(wire_d58_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905842(.data_in(wire_d58_41),.data_out(wire_d58_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905843(.data_in(wire_d58_42),.data_out(wire_d58_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905844(.data_in(wire_d58_43),.data_out(wire_d58_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905845(.data_in(wire_d58_44),.data_out(wire_d58_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905846(.data_in(wire_d58_45),.data_out(wire_d58_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905847(.data_in(wire_d58_46),.data_out(wire_d58_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905848(.data_in(wire_d58_47),.data_out(wire_d58_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905849(.data_in(wire_d58_48),.data_out(wire_d58_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905850(.data_in(wire_d58_49),.data_out(wire_d58_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905851(.data_in(wire_d58_50),.data_out(wire_d58_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905852(.data_in(wire_d58_51),.data_out(wire_d58_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905853(.data_in(wire_d58_52),.data_out(wire_d58_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905854(.data_in(wire_d58_53),.data_out(wire_d58_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905855(.data_in(wire_d58_54),.data_out(wire_d58_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905856(.data_in(wire_d58_55),.data_out(wire_d58_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905857(.data_in(wire_d58_56),.data_out(wire_d58_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905858(.data_in(wire_d58_57),.data_out(wire_d58_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905859(.data_in(wire_d58_58),.data_out(wire_d58_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905860(.data_in(wire_d58_59),.data_out(wire_d58_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905861(.data_in(wire_d58_60),.data_out(wire_d58_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905862(.data_in(wire_d58_61),.data_out(wire_d58_62),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905863(.data_in(wire_d58_62),.data_out(wire_d58_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905864(.data_in(wire_d58_63),.data_out(wire_d58_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905865(.data_in(wire_d58_64),.data_out(wire_d58_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905866(.data_in(wire_d58_65),.data_out(wire_d58_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905867(.data_in(wire_d58_66),.data_out(wire_d58_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905868(.data_in(wire_d58_67),.data_out(wire_d58_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905869(.data_in(wire_d58_68),.data_out(wire_d58_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905870(.data_in(wire_d58_69),.data_out(wire_d58_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905871(.data_in(wire_d58_70),.data_out(wire_d58_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905872(.data_in(wire_d58_71),.data_out(wire_d58_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905873(.data_in(wire_d58_72),.data_out(wire_d58_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905874(.data_in(wire_d58_73),.data_out(wire_d58_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905875(.data_in(wire_d58_74),.data_out(wire_d58_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905876(.data_in(wire_d58_75),.data_out(wire_d58_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905877(.data_in(wire_d58_76),.data_out(wire_d58_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905878(.data_in(wire_d58_77),.data_out(wire_d58_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905879(.data_in(wire_d58_78),.data_out(d_out58),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance600590(.data_in(d_in59),.data_out(wire_d59_0),.clk(clk),.rst(rst));            //channel 60
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance600591(.data_in(wire_d59_0),.data_out(wire_d59_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance600592(.data_in(wire_d59_1),.data_out(wire_d59_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance600593(.data_in(wire_d59_2),.data_out(wire_d59_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance600594(.data_in(wire_d59_3),.data_out(wire_d59_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance600595(.data_in(wire_d59_4),.data_out(wire_d59_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance600596(.data_in(wire_d59_5),.data_out(wire_d59_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance600597(.data_in(wire_d59_6),.data_out(wire_d59_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance600598(.data_in(wire_d59_7),.data_out(wire_d59_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance600599(.data_in(wire_d59_8),.data_out(wire_d59_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005910(.data_in(wire_d59_9),.data_out(wire_d59_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005911(.data_in(wire_d59_10),.data_out(wire_d59_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005912(.data_in(wire_d59_11),.data_out(wire_d59_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005913(.data_in(wire_d59_12),.data_out(wire_d59_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005914(.data_in(wire_d59_13),.data_out(wire_d59_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005915(.data_in(wire_d59_14),.data_out(wire_d59_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005916(.data_in(wire_d59_15),.data_out(wire_d59_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005917(.data_in(wire_d59_16),.data_out(wire_d59_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005918(.data_in(wire_d59_17),.data_out(wire_d59_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005919(.data_in(wire_d59_18),.data_out(wire_d59_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005920(.data_in(wire_d59_19),.data_out(wire_d59_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005921(.data_in(wire_d59_20),.data_out(wire_d59_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005922(.data_in(wire_d59_21),.data_out(wire_d59_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005923(.data_in(wire_d59_22),.data_out(wire_d59_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005924(.data_in(wire_d59_23),.data_out(wire_d59_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005925(.data_in(wire_d59_24),.data_out(wire_d59_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005926(.data_in(wire_d59_25),.data_out(wire_d59_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005927(.data_in(wire_d59_26),.data_out(wire_d59_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005928(.data_in(wire_d59_27),.data_out(wire_d59_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005929(.data_in(wire_d59_28),.data_out(wire_d59_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005930(.data_in(wire_d59_29),.data_out(wire_d59_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005931(.data_in(wire_d59_30),.data_out(wire_d59_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005932(.data_in(wire_d59_31),.data_out(wire_d59_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005933(.data_in(wire_d59_32),.data_out(wire_d59_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005934(.data_in(wire_d59_33),.data_out(wire_d59_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005935(.data_in(wire_d59_34),.data_out(wire_d59_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005936(.data_in(wire_d59_35),.data_out(wire_d59_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005937(.data_in(wire_d59_36),.data_out(wire_d59_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005938(.data_in(wire_d59_37),.data_out(wire_d59_38),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005939(.data_in(wire_d59_38),.data_out(wire_d59_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005940(.data_in(wire_d59_39),.data_out(wire_d59_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005941(.data_in(wire_d59_40),.data_out(wire_d59_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005942(.data_in(wire_d59_41),.data_out(wire_d59_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005943(.data_in(wire_d59_42),.data_out(wire_d59_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005944(.data_in(wire_d59_43),.data_out(wire_d59_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005945(.data_in(wire_d59_44),.data_out(wire_d59_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005946(.data_in(wire_d59_45),.data_out(wire_d59_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005947(.data_in(wire_d59_46),.data_out(wire_d59_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005948(.data_in(wire_d59_47),.data_out(wire_d59_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005949(.data_in(wire_d59_48),.data_out(wire_d59_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005950(.data_in(wire_d59_49),.data_out(wire_d59_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005951(.data_in(wire_d59_50),.data_out(wire_d59_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005952(.data_in(wire_d59_51),.data_out(wire_d59_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005953(.data_in(wire_d59_52),.data_out(wire_d59_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005954(.data_in(wire_d59_53),.data_out(wire_d59_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005955(.data_in(wire_d59_54),.data_out(wire_d59_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005956(.data_in(wire_d59_55),.data_out(wire_d59_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005957(.data_in(wire_d59_56),.data_out(wire_d59_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005958(.data_in(wire_d59_57),.data_out(wire_d59_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005959(.data_in(wire_d59_58),.data_out(wire_d59_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005960(.data_in(wire_d59_59),.data_out(wire_d59_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005961(.data_in(wire_d59_60),.data_out(wire_d59_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005962(.data_in(wire_d59_61),.data_out(wire_d59_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005963(.data_in(wire_d59_62),.data_out(wire_d59_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005964(.data_in(wire_d59_63),.data_out(wire_d59_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005965(.data_in(wire_d59_64),.data_out(wire_d59_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005966(.data_in(wire_d59_65),.data_out(wire_d59_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005967(.data_in(wire_d59_66),.data_out(wire_d59_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005968(.data_in(wire_d59_67),.data_out(wire_d59_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005969(.data_in(wire_d59_68),.data_out(wire_d59_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005970(.data_in(wire_d59_69),.data_out(wire_d59_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005971(.data_in(wire_d59_70),.data_out(wire_d59_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005972(.data_in(wire_d59_71),.data_out(wire_d59_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005973(.data_in(wire_d59_72),.data_out(wire_d59_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005974(.data_in(wire_d59_73),.data_out(wire_d59_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005975(.data_in(wire_d59_74),.data_out(wire_d59_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005976(.data_in(wire_d59_75),.data_out(wire_d59_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005977(.data_in(wire_d59_76),.data_out(wire_d59_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005978(.data_in(wire_d59_77),.data_out(wire_d59_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005979(.data_in(wire_d59_78),.data_out(d_out59),.clk(clk),.rst(rst));


endmodule