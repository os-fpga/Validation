module BUF_X1(A, Y);
input A;
output Y;
assign Y = A;
endmodule